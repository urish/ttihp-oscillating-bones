* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] VAPWR VDPWR VGND
X0 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t20 VGND.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X1 VAPWR.t41 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VAPWR.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X2 VAPWR.t15 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VAPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X3 a_13289_43697# uo_out[2].t2 VDPWR.t59 VDPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X4 a_16868_43697# a_17160_43997# a_17111_44089# VDPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X5 a_16596_43697# a_16868_43697# VGND.t63 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VDPWR.t41 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND.t60 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X8 a_15221_43697# uo_out[1].t2 VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9 VDPWR.t65 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VDPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X10 a_15179_44089# a_14664_43697# VDPWR.t71 VDPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VGND.t5 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_6.A VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X12 a_17360_43697# a_17160_43997# a_17509_43723# VGND.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X13 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VAPWR.t25 VAPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X14 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VAPWR.t3 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X15 a_15577_43723# a_15357_43723# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X16 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VAPWR.t5 VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X17 VGND.t86 a_14664_43697# uo_out[2].t0 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X18 VDPWR.t25 a_13289_43697# a_13296_43997# VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X19 VGND.t80 a_15221_43697# a_15228_43997# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VAPWR.t11 VAPWR.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X21 a_13843_43723# a_13296_43997# a_13496_43697# VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X22 a_16501_43697# a_16596_43697# VGND.t26 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X23 a_12637_43697# a_12732_43697# VDPWR.t39 VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X24 a_17289_43723# a_17153_43697# a_16868_43697# VDPWR.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X25 a_13224_43723# a_12732_43697# VGND.t55 VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 VGND.t62 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VGND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X27 VGND.t48 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X28 VDPWR.t69 a_14664_43697# uo_out[2].t1 VDPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X29 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VAPWR.t13 VAPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X30 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t35 VGND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X31 a_15156_43723# a_14664_43697# VGND.t85 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X32 a_17707_43723# a_17153_43697# a_17360_43697# VGND.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X33 a_14936_43697# a_15228_43997# a_15179_44089# VDPWR.t5 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X34 a_13289_43697# uo_out[2].t3 VGND.t31 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X35 VGND.t79 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X36 a_14664_43697# a_14936_43697# VGND.t44 VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X37 VGND.t57 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X38 VGND.t3 a_13496_43697# a_13425_43723# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X39 VAPWR.t17 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VAPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X40 uo_out[0].t1 skullfet_level_shifter.A VGND.t69 VGND.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X41 a_13247_44089# a_12732_43697# VDPWR.t37 VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X42 a_15221_43697# uo_out[1].t3 VGND.t16 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 a_15428_43697# a_15228_43997# a_15577_43723# VGND.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X44 VGND.t28 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X45 a_13645_43723# a_13425_43723# VGND.t42 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X46 VGND.t39 a_15428_43697# a_15357_43723# VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X47 VGND.t53 a_12732_43697# uo_out[3].t1 VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X48 VDPWR.t43 a_17360_43697# a_17289_43723# VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X49 a_16868_43697# a_17153_43697# a_17088_43723# VGND.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X50 a_14664_43697# a_14936_43697# VDPWR.t31 VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X51 VAPWR.t9 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VAPWR.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X52 VGND.t41 a_13289_43697# a_13296_43997# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X53 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_8.A VAPWR.t33 VAPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X54 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VAPWR.t35 VAPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X55 a_14569_43697# a_14664_43697# VGND.t84 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X56 a_15604_44089# a_15357_43723# VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X57 a_15357_43723# a_15221_43697# a_14936_43697# VDPWR.t63 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X58 a_15428_43697# a_15221_43697# a_15604_44089# VDPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X59 a_12732_43697# a_13004_43697# VGND.t73 VGND.t72 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X60 VGND.t12 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X61 VDPWR.t57 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VDPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X62 VDPWR.t35 a_12732_43697# uo_out[3].t0 VDPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X63 a_17289_43723# a_17160_43997# a_16868_43697# VGND.t15 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X64 a_17153_43697# uo_out[0].t2 VDPWR.t73 VDPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X65 a_17536_44089# a_17289_43723# VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X66 VGND.t22 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X67 a_17360_43697# a_17153_43697# a_17536_44089# VDPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X68 a_17111_44089# a_16596_43697# VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X69 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VAPWR.t27 VAPWR.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X70 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VAPWR.t37 VAPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X71 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t30 VGND.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X72 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VAPWR.t29 VAPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X73 a_15775_43723# a_15221_43697# a_15428_43697# VGND.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X74 a_13004_43697# a_13296_43997# a_13247_44089# VDPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X75 VDPWR.t33 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X76 VGND.t71 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_9.A VGND.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X77 a_12732_43697# a_13004_43697# VDPWR.t53 VDPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X78 VGND.t75 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X79 VGND.t76 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X80 a_16501_43697# a_16596_43697# VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X81 a_13496_43697# a_13296_43997# a_13645_43723# VGND.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X82 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_4.A VAPWR.t23 VAPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X83 ring_0/skullfet_inverter_8.A skullfet_level_shifter.A VAPWR.t31 VAPWR.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X84 VGND.t78 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X85 VDPWR.t21 a_15428_43697# a_15357_43723# VDPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X86 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t37 VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X87 VDPWR.t11 a_17153_43697# a_17160_43997# VDPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X88 VGND.t65 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X89 a_14936_43697# a_15221_43697# a_15156_43723# VGND.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X90 VDPWR.t51 skullfet_level_shifter.A uo_out[0].t0 VDPWR.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X91 VGND.t7 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X92 a_12637_43697# a_12732_43697# VGND.t51 VGND.t50 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X93 VGND.t83 ring_0/skullfet_inverter_6.A skullfet_level_shifter.A VGND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X94 a_13672_44089# a_13425_43723# VDPWR.t29 VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X95 a_13425_43723# a_13296_43997# a_13004_43697# VGND.t13 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X96 VGND.t18 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X97 a_13425_43723# a_13289_43697# a_13004_43697# VDPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X98 a_13496_43697# a_13289_43697# a_13672_44089# VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X99 VDPWR.t45 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X100 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t33 VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X101 VGND.t46 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_5.A VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X102 VDPWR.t55 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VDPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X103 VGND.t67 skullfet_level_shifter.A ring_0/skullfet_inverter_8.A VGND.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X104 a_15357_43723# a_15228_43997# a_14936_43697# VGND.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X105 a_17153_43697# uo_out[0].t3 VGND.t87 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X106 VAPWR.t21 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VAPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X107 a_17509_43723# a_17289_43723# VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X108 VGND.t25 a_16596_43697# uo_out[1].t1 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X109 a_13843_43723# a_13289_43697# a_13496_43697# VGND.t8 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X110 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t89 VGND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X111 VGND.t59 a_17360_43697# a_17289_43723# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X112 VGND.t49 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X113 VDPWR.t61 a_15221_43697# a_15228_43997# VDPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X114 VGND.t81 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X115 VAPWR.t19 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VAPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X116 a_15775_43723# a_15228_43997# a_15428_43697# VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X117 a_13004_43697# a_13289_43697# a_13224_43723# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X118 skullfet_level_shifter.A ring_0/skullfet_inverter_6.A VAPWR.t39 VAPWR.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X119 a_16596_43697# a_16868_43697# VDPWR.t47 VDPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X120 a_14569_43697# a_14664_43697# VDPWR.t67 VDPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X121 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VAPWR.t7 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X122 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_5.A VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X123 a_17707_43723# a_17160_43997# a_17360_43697# VDPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X124 VDPWR.t15 a_16596_43697# uo_out[1].t0 VDPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X125 VDPWR.t3 a_13496_43697# a_13425_43723# VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X126 VGND.t14 a_17153_43697# a_17160_43997# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X127 a_17088_43723# a_16596_43697# VGND.t23 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 VGND.n425 VGND.n424 570379
R1 VGND.n130 VGND.n129 570263
R2 VGND.n129 VGND.n3 194461
R3 VGND.n425 VGND.n24 194343
R4 VGND.n130 VGND.n78 192789
R5 VGND.n424 VGND.n423 192674
R6 VGND.n158 VGND.n156 57198.5
R7 VGND.n132 VGND.n131 54022.2
R8 VGND.n26 VGND.n25 54013.8
R9 VGND.n472 VGND.n4 36049.1
R10 VGND.n423 VGND.t82 32282.1
R11 VGND.n102 VGND.n78 30458.6
R12 VGND.n77 VGND.n3 30455.9
R13 VGND.n325 VGND.n24 30451.1
R14 VGND.n423 VGND.n26 30163.7
R15 VGND.n99 VGND.n78 30163.7
R16 VGND.n137 VGND.n75 27183.9
R17 VGND.t11 VGND.n152 22572.7
R18 VGND.n152 VGND.n151 19011.9
R19 VGND.n322 VGND.t15 16545.7
R20 VGND.t56 VGND.n158 14642.2
R21 VGND.n136 VGND.n132 14211.6
R22 VGND.n334 VGND.n156 13525.9
R23 VGND.n424 VGND.n25 13282
R24 VGND.n131 VGND.n130 13281.9
R25 VGND.n135 VGND.n74 12582
R26 VGND.n472 VGND.n471 11835.1
R27 VGND.n322 VGND.n321 11079.9
R28 VGND.n138 VGND.n74 8411.7
R29 VGND.n138 VGND.n137 7811.4
R30 VGND.n325 VGND.n25 6174.02
R31 VGND.n131 VGND.n77 6169.66
R32 VGND.n322 VGND.n318 5759.37
R33 VGND.n471 VGND.t27 5611.54
R34 VGND.n140 VGND.n68 5579.62
R35 VGND.n132 VGND.n74 5351.68
R36 VGND.n135 VGND.n134 4937.85
R37 VGND.n140 VGND.n139 4845.05
R38 VGND.n69 VGND.n7 4441.64
R39 VGND.n334 VGND.n325 4412.94
R40 VGND.n334 VGND.n157 4224.13
R41 VGND.n136 VGND.n135 3889.67
R42 VGND.t68 VGND.n27 3753.63
R43 VGND.n128 VGND.n3 3692.64
R44 VGND.n77 VGND.n75 3402.31
R45 VGND.n471 VGND.n470 3172.32
R46 VGND.n469 VGND.t17 2863.06
R47 VGND.n422 VGND.n421 2777.19
R48 VGND.n422 VGND.n27 2407.29
R49 VGND.n322 VGND 2376.85
R50 VGND.n426 VGND.n24 2322.17
R51 VGND.t64 VGND.n8 2286.05
R52 VGND.t36 VGND.n472 2076.87
R53 VGND.n71 VGND.n70 2060.84
R54 VGND.n333 VGND.n331 1852.32
R55 VGND.n334 VGND.n324 1851.9
R56 VGND.n7 VGND.n6 1798.88
R57 VGND.n322 VGND.n27 1764.6
R58 VGND.n470 VGND.n7 1655.02
R59 VGND.n332 VGND.n9 1554.7
R60 VGND.n139 VGND.n138 1540.61
R61 VGND.n134 VGND.t29 1523.34
R62 VGND.n151 VGND.t21 1449.81
R63 VGND.n155 VGND.n154 1403.85
R64 VGND.n72 VGND.n71 1385.1
R65 VGND.n321 VGND.t4 1309.34
R66 VGND.n139 VGND.t21 1230.65
R67 VGND.n137 VGND.n136 1226.09
R68 VGND.t74 VGND.n68 1163.46
R69 VGND.t29 VGND.n132 1127.76
R70 VGND.n129 VGND.t88 1089.82
R71 VGND.t66 VGND.n425 1089.82
R72 VGND.n132 VGND.n76 954.316
R73 VGND.n340 VGND.n26 938.943
R74 VGND.n6 VGND.t27 898.419
R75 VGND.t54 VGND.t72 809.293
R76 VGND.t32 VGND.n3 807.455
R77 VGND.t52 VGND.t50 800.774
R78 VGND.n102 VGND.t34 771.376
R79 VGND.n157 VGND.n26 769.477
R80 VGND.n273 VGND.n24 722.872
R81 VGND.n155 VGND.n68 712.85
R82 VGND.n99 VGND.t19 711.236
R83 VGND.t6 VGND.n155 710.678
R84 VGND.t45 VGND.n26 710.202
R85 VGND.n333 VGND.n332 641.15
R86 VGND.n158 VGND.n24 604.66
R87 VGND.n154 VGND.t11 599.504
R88 VGND.n317 VGND.n159 595.942
R89 VGND.n317 VGND.n316 595.942
R90 VGND.n328 VGND.n327 585
R91 VGND.n330 VGND.n329 585
R92 VGND.n466 VGND.n465 585
R93 VGND.n469 VGND.n468 585
R94 VGND.n6 VGND.n5 585
R95 VGND.n474 VGND.n473 585
R96 VGND.n128 VGND.n127 585
R97 VGND.n101 VGND.n100 585
R98 VGND.n96 VGND.n76 585
R99 VGND.n104 VGND.n103 585
R100 VGND.n142 VGND.n141 585
R101 VGND.n321 VGND.n320 585
R102 VGND.n427 VGND.n426 585
R103 VGND.n274 VGND.n273 585
R104 VGND.n324 VGND.n323 585
R105 VGND.n336 VGND.n335 585
R106 VGND.n154 VGND.n153 585
R107 VGND.n145 VGND.n144 585
R108 VGND.n151 VGND.n150 585
R109 VGND.n134 VGND.n133 585
R110 VGND.n103 VGND.n102 580.986
R111 VGND.n27 VGND.n24 561.288
R112 VGND.n71 VGND.n7 558.698
R113 VGND.n144 VGND.t74 546.268
R114 VGND.n101 VGND.n99 541.24
R115 VGND.n273 VGND.t68 459.25
R116 VGND.t13 VGND.t40 451.5
R117 VGND.n152 VGND.n69 435.567
R118 VGND.n152 VGND.t61 433.632
R119 VGND.t2 VGND.t13 430.204
R120 VGND.t82 VGND.n422 424.454
R121 VGND.n152 VGND.n8 416.322
R122 VGND.n70 VGND.n69 416.322
R123 VGND.t40 VGND.t54 404.647
R124 VGND.t50 VGND.t56 404.647
R125 VGND.n318 VGND.t2 370.572
R126 VGND.t72 VGND.t52 357.793
R127 VGND.n334 VGND.n333 343.485
R128 VGND.n318 VGND 343.437
R129 VGND.t64 VGND.n469 340.748
R130 VGND.n157 VGND.t47 338.3
R131 VGND.n142 VGND.t61 332.805
R132 VGND.t21 VGND.n70 330.817
R133 VGND.n331 VGND.n328 308.387
R134 VGND.t88 VGND.n128 304.548
R135 VGND.n426 VGND.t66 304.548
R136 VGND.n332 VGND.n8 294.779
R137 VGND.n323 VGND.t46 282.13
R138 VGND.n336 VGND.t7 282.13
R139 VGND.n145 VGND.t75 282.13
R140 VGND.n427 VGND.t67 282.13
R141 VGND.n329 VGND.t78 282.13
R142 VGND.n468 VGND.t65 282.13
R143 VGND.n327 VGND.t71 282.13
R144 VGND.n340 VGND.t48 282.13
R145 VGND.n320 VGND.t5 282.13
R146 VGND.n421 VGND.t83 282.13
R147 VGND.n274 VGND.t69 281.841
R148 VGND.n153 VGND.t12 281.839
R149 VGND.n150 VGND.t22 281.839
R150 VGND.n104 VGND.t33 281.839
R151 VGND.n465 VGND.t18 281.839
R152 VGND.n5 VGND.t28 281.839
R153 VGND.n474 VGND.t37 281.839
R154 VGND.n127 VGND.t89 281.839
R155 VGND.n96 VGND.t20 281.839
R156 VGND.n100 VGND.t35 281.839
R157 VGND.n133 VGND.t30 281.839
R158 VGND.n141 VGND.t62 281.839
R159 VGND.n144 VGND.n143 259.74
R160 VGND.n238 VGND.t85 251
R161 VGND.n205 VGND.t23 251
R162 VGND.n296 VGND.t55 251
R163 VGND.n225 VGND.t76 243.028
R164 VGND.n192 VGND.t79 243.028
R165 VGND.n309 VGND.t81 243.028
R166 VGND.n334 VGND.n322 222.743
R167 VGND.n143 VGND.n140 221.165
R168 VGND.n240 VGND.n165 218.506
R169 VGND.n179 VGND.n178 218.506
R170 VGND.n261 VGND.n260 218.506
R171 VGND.n246 VGND.n162 200.201
R172 VGND.n176 VGND.n175 200.201
R173 VGND.n264 VGND.n263 200.201
R174 VGND.n174 VGND.n173 199.739
R175 VGND.n188 VGND.n187 199.739
R176 VGND.n252 VGND.n251 199.739
R177 VGND.n231 VGND.n169 199.53
R178 VGND.n198 VGND.n183 199.53
R179 VGND.n303 VGND.n256 199.53
R180 VGND.n75 VGND.n4 194.254
R181 VGND.t34 VGND.n101 194.014
R182 VGND.n324 VGND.t45 192.522
R183 VGND.n103 VGND.t32 188.929
R184 VGND.t19 VGND.n76 179.65
R185 VGND.t70 VGND.n24 178.903
R186 VGND.n331 VGND.t77 147.839
R187 VGND.n330 VGND.n9 142.013
R188 VGND.n473 VGND.t36 140.379
R189 VGND.n328 VGND.t70 137.305
R190 VGND.n335 VGND.t6 124.846
R191 VGND VGND.t8 119.269
R192 VGND.t77 VGND.n330 113.463
R193 VGND.t9 VGND.n156 96.261
R194 VGND.t17 VGND.n466 94.4922
R195 VGND.t21 VGND.n72 85.506
R196 VGND.t9 VGND.t58 83.7375
R197 VGND.n169 VGND.t39 74.8666
R198 VGND.n183 VGND.t59 74.8666
R199 VGND.n256 VGND.t3 74.8666
R200 VGND.n470 VGND.t64 67.3773
R201 VGND.n162 VGND.t84 54.2862
R202 VGND.n175 VGND.t26 54.2862
R203 VGND.n263 VGND.t51 54.2862
R204 VGND VGND.t9 49.8097
R205 VGND.n473 VGND.n3 46.3668
R206 VGND.n335 VGND.n334 41.2363
R207 VGND.n169 VGND.t1 40.0005
R208 VGND.n183 VGND.t10 40.0005
R209 VGND.n256 VGND.t42 40.0005
R210 VGND.n173 VGND.t16 38.5719
R211 VGND.n173 VGND.t80 38.5719
R212 VGND.n187 VGND.t87 38.5719
R213 VGND.n187 VGND.t14 38.5719
R214 VGND.n251 VGND.t31 38.5719
R215 VGND.n251 VGND.t41 38.5719
R216 VGND.n241 VGND.n163 34.6358
R217 VGND.n245 VGND.n163 34.6358
R218 VGND.n233 VGND.n232 34.6358
R219 VGND.n233 VGND.n167 34.6358
R220 VGND.n237 VGND.n167 34.6358
R221 VGND.n226 VGND.n171 34.6358
R222 VGND.n230 VGND.n171 34.6358
R223 VGND.n210 VGND.n209 34.6358
R224 VGND.n211 VGND.n210 34.6358
R225 VGND.n200 VGND.n199 34.6358
R226 VGND.n200 VGND.n181 34.6358
R227 VGND.n204 VGND.n181 34.6358
R228 VGND.n193 VGND.n185 34.6358
R229 VGND.n197 VGND.n185 34.6358
R230 VGND.n308 VGND.n254 34.6358
R231 VGND.n304 VGND.n254 34.6358
R232 VGND.n302 VGND.n257 34.6358
R233 VGND.n298 VGND.n257 34.6358
R234 VGND.n298 VGND.n297 34.6358
R235 VGND.n292 VGND.n291 34.6358
R236 VGND.n291 VGND.n290 34.6358
R237 VGND.n240 VGND.n239 32.7534
R238 VGND.n206 VGND.n179 32.7534
R239 VGND.n295 VGND.n261 32.7534
R240 VGND.t0 VGND.t38 31.6138
R241 VGND.n239 VGND.n238 31.2476
R242 VGND.n206 VGND.n205 31.2476
R243 VGND.n296 VGND.n295 31.2476
R244 VGND.n466 VGND.n9 31.2108
R245 VGND.n231 VGND.n230 30.8711
R246 VGND.n198 VGND.n197 30.8711
R247 VGND.n304 VGND.n303 30.8711
R248 VGND.n226 VGND.n225 27.4829
R249 VGND.n193 VGND.n192 27.4829
R250 VGND.n309 VGND.n308 27.4829
R251 VGND.n162 VGND.t60 25.9346
R252 VGND.n175 VGND.t49 25.9346
R253 VGND.n263 VGND.t57 25.9346
R254 VGND.n165 VGND.t44 24.9236
R255 VGND.n165 VGND.t86 24.9236
R256 VGND.n178 VGND.t63 24.9236
R257 VGND.n178 VGND.t25 24.9236
R258 VGND.n260 VGND.t73 24.9236
R259 VGND.n260 VGND.t53 24.9236
R260 VGND.n247 VGND.n160 23.7181
R261 VGND.n246 VGND.n245 23.7181
R262 VGND.n220 VGND.n219 23.7181
R263 VGND.n216 VGND.n215 23.7181
R264 VGND.n211 VGND.n176 23.7181
R265 VGND.n315 VGND.n314 23.7181
R266 VGND.n290 VGND.n264 23.7181
R267 VGND.n143 VGND.n142 23.5015
R268 VGND.t43 VGND.n317 22.992
R269 VGND.n224 VGND.n174 22.9652
R270 VGND.n225 VGND.n224 22.9652
R271 VGND.n191 VGND.n188 22.9652
R272 VGND.n192 VGND.n191 22.9652
R273 VGND.n310 VGND.n252 22.9652
R274 VGND.n310 VGND.n309 22.9652
R275 VGND.t9 VGND.t15 22.8379
R276 VGND.n238 VGND.n237 22.2123
R277 VGND.n205 VGND.n204 22.2123
R278 VGND.n297 VGND.n296 22.2123
R279 VGND.n72 VGND.n4 21.5982
R280 VGND.n247 VGND.n246 21.4593
R281 VGND.n220 VGND.n174 21.4593
R282 VGND.n215 VGND.n176 21.4593
R283 VGND.n314 VGND.n252 21.4593
R284 VGND.n149 VGND.n73 21.2541
R285 VGND.n476 VGND.n475 16.3975
R286 VGND.n323 VGND.n48 13.2958
R287 VGND.n337 VGND.n336 13.2958
R288 VGND.n146 VGND.n145 13.2958
R289 VGND.n428 VGND.n427 13.2958
R290 VGND.n329 VGND.n10 13.2958
R291 VGND.n468 VGND.n467 13.2958
R292 VGND.n327 VGND.n326 13.2958
R293 VGND.n341 VGND.n340 13.2958
R294 VGND.n320 VGND.n319 13.2958
R295 VGND.n421 VGND.n420 13.2958
R296 VGND VGND.n274 13.2396
R297 VGND.n153 VGND 13.2396
R298 VGND.n150 VGND 13.2396
R299 VGND.n465 VGND 13.2396
R300 VGND.n5 VGND 13.2396
R301 VGND VGND.n474 13.2396
R302 VGND.n127 VGND 13.2396
R303 VGND VGND.n96 13.2396
R304 VGND.n100 VGND 13.2396
R305 VGND VGND.n104 13.2396
R306 VGND.n133 VGND 13.2396
R307 VGND.n141 VGND 13.2396
R308 VGND.n283 VGND 12.8296
R309 VGND VGND.n287 11.784
R310 VGND.n232 VGND.n231 10.5417
R311 VGND.n199 VGND.n198 10.5417
R312 VGND.n303 VGND.n302 10.5417
R313 VGND.n476 VGND 9.61512
R314 VGND.n290 VGND.n289 9.3005
R315 VGND.n291 VGND.n262 9.3005
R316 VGND.n293 VGND.n292 9.3005
R317 VGND.n295 VGND.n294 9.3005
R318 VGND.n296 VGND.n259 9.3005
R319 VGND.n297 VGND.n258 9.3005
R320 VGND.n299 VGND.n298 9.3005
R321 VGND.n300 VGND.n257 9.3005
R322 VGND.n302 VGND.n301 9.3005
R323 VGND.n303 VGND.n255 9.3005
R324 VGND.n305 VGND.n304 9.3005
R325 VGND.n306 VGND.n254 9.3005
R326 VGND.n308 VGND.n307 9.3005
R327 VGND.n309 VGND.n253 9.3005
R328 VGND.n311 VGND.n310 9.3005
R329 VGND.n312 VGND.n252 9.3005
R330 VGND.n314 VGND.n313 9.3005
R331 VGND.n315 VGND.n250 9.3005
R332 VGND.n191 VGND.n190 9.3005
R333 VGND.n192 VGND.n186 9.3005
R334 VGND.n194 VGND.n193 9.3005
R335 VGND.n195 VGND.n185 9.3005
R336 VGND.n197 VGND.n196 9.3005
R337 VGND.n198 VGND.n184 9.3005
R338 VGND.n199 VGND.n182 9.3005
R339 VGND.n201 VGND.n200 9.3005
R340 VGND.n202 VGND.n181 9.3005
R341 VGND.n204 VGND.n203 9.3005
R342 VGND.n205 VGND.n180 9.3005
R343 VGND.n207 VGND.n206 9.3005
R344 VGND.n209 VGND.n208 9.3005
R345 VGND.n210 VGND.n177 9.3005
R346 VGND.n212 VGND.n211 9.3005
R347 VGND.n213 VGND.n176 9.3005
R348 VGND.n215 VGND.n214 9.3005
R349 VGND.n217 VGND.n216 9.3005
R350 VGND.n219 VGND.n218 9.3005
R351 VGND.n221 VGND.n220 9.3005
R352 VGND.n222 VGND.n174 9.3005
R353 VGND.n224 VGND.n223 9.3005
R354 VGND.n225 VGND.n172 9.3005
R355 VGND.n227 VGND.n226 9.3005
R356 VGND.n228 VGND.n171 9.3005
R357 VGND.n230 VGND.n229 9.3005
R358 VGND.n231 VGND.n170 9.3005
R359 VGND.n232 VGND.n168 9.3005
R360 VGND.n234 VGND.n233 9.3005
R361 VGND.n235 VGND.n167 9.3005
R362 VGND.n237 VGND.n236 9.3005
R363 VGND.n238 VGND.n166 9.3005
R364 VGND.n239 VGND.n164 9.3005
R365 VGND.n242 VGND.n241 9.3005
R366 VGND.n243 VGND.n163 9.3005
R367 VGND.n245 VGND.n244 9.3005
R368 VGND.n246 VGND.n161 9.3005
R369 VGND.n248 VGND.n247 9.3005
R370 VGND.n249 VGND.n160 9.3005
R371 VGND.n463 VGND.n462 9.1888
R372 VGND VGND.n149 9.01182
R373 VGND.n339 VGND.n338 8.65869
R374 VGND.t8 VGND.t0 8.62232
R375 VGND.n147 VGND.n146 8.4976
R376 VGND VGND.n464 8.23872
R377 VGND.n148 VGND 8.06793
R378 VGND.n338 VGND.n337 7.59474
R379 VGND.n467 VGND.n1 7.53106
R380 VGND.n189 VGND.n188 7.12576
R381 VGND.n288 VGND.n264 7.12063
R382 VGND.n475 VGND 7.08005
R383 VGND VGND.n67 6.79835
R384 VGND.n463 VGND.n10 6.59477
R385 VGND.n342 VGND.n341 6.49817
R386 VGND.n216 VGND.n159 6.367
R387 VGND.n316 VGND.n315 6.367
R388 VGND.n316 VGND.n160 6.367
R389 VGND.n219 VGND.n159 6.367
R390 VGND VGND.n73 6.28926
R391 VGND VGND.n126 6.23801
R392 VGND.n326 VGND.n11 6.09911
R393 VGND.n361 VGND.n48 6.00714
R394 VGND VGND.n98 5.93135
R395 VGND.n97 VGND 5.83554
R396 VGND.n420 VGND.n419 5.80344
R397 VGND.n105 VGND 5.75987
R398 VGND.n319 VGND.n28 5.70397
R399 VGND.n429 VGND.n428 5.56083
R400 VGND.n275 VGND.n0 4.70536
R401 VGND.t58 VGND.t24 3.80673
R402 VGND.n0 VGND 3.44325
R403 VGND.n97 VGND.n73 3.41091
R404 VGND.n479 VGND 3.36335
R405 VGND.n338 VGND.n67 2.9742
R406 VGND VGND.n479 2.3855
R407 VGND.n464 VGND.n463 2.0669
R408 VGND.n241 VGND.n240 1.88285
R409 VGND.n209 VGND.n179 1.88285
R410 VGND.n292 VGND.n261 1.88285
R411 VGND.t38 VGND.t43 1.43747
R412 VGND.n149 VGND.n148 1.34683
R413 VGND.n98 VGND.n97 1.13252
R414 VGND.n464 VGND.n1 1.02753
R415 VGND.n148 VGND.n147 0.99238
R416 VGND.n147 VGND.n67 0.965475
R417 VGND.n381 VGND.n28 0.8755
R418 VGND.n475 VGND.n2 0.827423
R419 VGND.n477 VGND.n476 0.715835
R420 VGND.n106 VGND.n98 0.576786
R421 VGND.n478 VGND.n477 0.520466
R422 VGND.n384 VGND.n383 0.454101
R423 VGND.n265 uo_out[4] 0.39812
R424 VGND.n265 uo_out[5] 0.2684
R425 VGND.n266 uo_out[6] 0.2684
R426 VGND.n267 uo_out[7] 0.2684
R427 VGND.n268 uio_out[0] 0.2684
R428 VGND.n269 uio_out[1] 0.2684
R429 VGND.n270 uio_out[2] 0.2684
R430 VGND.n271 uio_out[3] 0.2684
R431 VGND.n272 uio_out[4] 0.2684
R432 VGND.n286 uio_out[5] 0.2684
R433 VGND.n285 uio_out[6] 0.2684
R434 VGND.n284 uio_out[7] 0.2684
R435 VGND.n282 uio_oe[0] 0.2684
R436 VGND.n281 uio_oe[1] 0.2684
R437 VGND.n280 uio_oe[2] 0.2684
R438 VGND.n279 uio_oe[3] 0.2684
R439 VGND.n278 uio_oe[4] 0.2684
R440 VGND.n277 uio_oe[5] 0.2684
R441 VGND.n276 uio_oe[6] 0.2684
R442 VGND.n275 uio_oe[7] 0.2684
R443 VGND.n381 VGND.n380 0.240762
R444 VGND.n380 VGND.n379 0.212286
R445 VGND.n123 VGND.n79 0.173819
R446 VGND.n379 VGND.n378 0.17131
R447 VGND.n107 VGND.n106 0.167466
R448 VGND.n462 VGND.n461 0.160547
R449 VGND.n288 VGND 0.152603
R450 VGND.n378 VGND.n377 0.15242
R451 VGND.n289 VGND.n288 0.148519
R452 VGND.n124 VGND.n2 0.14598
R453 VGND.n190 VGND.n189 0.143396
R454 VGND.n377 VGND.n376 0.137604
R455 VGND.n382 VGND.n381 0.135859
R456 VGND.n380 VGND.n29 0.135168
R457 VGND.n378 VGND.n31 0.134528
R458 VGND.n383 VGND.n28 0.13451
R459 VGND.n379 VGND.n30 0.134478
R460 VGND.n376 VGND.n33 0.133139
R461 VGND.n377 VGND.n32 0.133097
R462 VGND.n374 VGND.n35 0.131785
R463 VGND.n375 VGND.n34 0.13175
R464 VGND.n371 VGND.n38 0.130416
R465 VGND.n372 VGND.n37 0.130388
R466 VGND.n373 VGND.n36 0.130361
R467 VGND.n266 VGND.n265 0.13022
R468 VGND.n267 VGND.n266 0.13022
R469 VGND.n268 VGND.n267 0.13022
R470 VGND.n269 VGND.n268 0.13022
R471 VGND.n270 VGND.n269 0.13022
R472 VGND.n271 VGND.n270 0.13022
R473 VGND.n272 VGND.n271 0.13022
R474 VGND.n286 VGND.n285 0.13022
R475 VGND.n285 VGND.n284 0.13022
R476 VGND.n282 VGND.n281 0.13022
R477 VGND.n281 VGND.n280 0.13022
R478 VGND.n280 VGND.n279 0.13022
R479 VGND.n279 VGND.n278 0.13022
R480 VGND.n278 VGND.n277 0.13022
R481 VGND.n277 VGND.n276 0.13022
R482 VGND.n276 VGND.n275 0.13022
R483 VGND.n107 VGND.n95 0.129737
R484 VGND.n109 VGND.n93 0.129051
R485 VGND.n108 VGND.n94 0.129031
R486 VGND.n368 VGND.n41 0.129031
R487 VGND.n369 VGND.n40 0.129011
R488 VGND.n370 VGND.n39 0.128992
R489 VGND.n367 VGND.n42 0.128325
R490 VGND.n112 VGND.n90 0.127655
R491 VGND.n111 VGND.n91 0.127643
R492 VGND.n110 VGND.n92 0.127631
R493 VGND.n461 VGND.n460 0.127299
R494 VGND.n459 VGND.n12 0.127286
R495 VGND.n458 VGND.n457 0.127273
R496 VGND.n115 VGND.n87 0.126953
R497 VGND.n114 VGND.n88 0.126945
R498 VGND.n113 VGND.n89 0.126937
R499 VGND.n417 VGND.n386 0.12692
R500 VGND.n365 VGND.n44 0.12692
R501 VGND.n418 VGND.n385 0.126912
R502 VGND.n366 VGND.n43 0.126912
R503 VGND.n456 VGND.n13 0.126374
R504 VGND.n453 VGND.n14 0.126362
R505 VGND.n120 VGND.n82 0.126244
R506 VGND.n118 VGND.n84 0.126235
R507 VGND.n117 VGND.n85 0.126231
R508 VGND.n116 VGND.n86 0.126227
R509 VGND.n414 VGND.n389 0.126218
R510 VGND.n362 VGND.n47 0.126218
R511 VGND.n415 VGND.n388 0.126214
R512 VGND.n363 VGND.n46 0.126214
R513 VGND.n416 VGND.n387 0.12621
R514 VGND.n364 VGND.n45 0.12621
R515 VGND.n376 VGND.n375 0.126068
R516 VGND.n413 VGND.n390 0.1255
R517 VGND.n412 VGND.n391 0.1255
R518 VGND.n411 VGND.n392 0.1255
R519 VGND.n449 VGND.n448 0.1255
R520 VGND.n452 VGND.n451 0.1255
R521 VGND.n455 VGND.n454 0.1255
R522 VGND.n122 VGND.n80 0.1255
R523 VGND.n358 VGND.n51 0.1255
R524 VGND.n359 VGND.n50 0.1255
R525 VGND.n360 VGND.n49 0.1255
R526 VGND.n410 VGND.n393 0.124773
R527 VGND.n357 VGND.n52 0.124773
R528 VGND.n408 VGND.n395 0.124765
R529 VGND.n119 VGND.n83 0.124765
R530 VGND.n355 VGND.n54 0.124765
R531 VGND.n406 VGND.n397 0.124756
R532 VGND.n121 VGND.n81 0.124756
R533 VGND.n353 VGND.n56 0.124756
R534 VGND.n409 VGND.n394 0.124038
R535 VGND.n356 VGND.n53 0.124038
R536 VGND.n441 VGND.n18 0.123887
R537 VGND.n444 VGND.n17 0.123866
R538 VGND.n447 VGND.n16 0.123844
R539 VGND.n450 VGND.n15 0.123822
R540 VGND.n124 VGND.n123 0.123412
R541 VGND.n407 VGND.n396 0.123294
R542 VGND.n354 VGND.n55 0.123294
R543 VGND.n405 VGND.n398 0.123268
R544 VGND.n352 VGND.n57 0.123268
R545 VGND.n404 VGND.n399 0.123254
R546 VGND.n351 VGND.n58 0.123254
R547 VGND.n403 VGND.n400 0.123241
R548 VGND.n350 VGND.n59 0.123241
R549 VGND.n23 VGND.n22 0.123213
R550 VGND.n348 VGND.n61 0.123213
R551 VGND.n431 VGND.n430 0.123199
R552 VGND.n347 VGND.n62 0.123199
R553 VGND.n432 VGND.n21 0.123185
R554 VGND.n346 VGND.n63 0.123185
R555 VGND.n434 VGND.n433 0.123171
R556 VGND.n345 VGND.n64 0.123171
R557 VGND.n437 VGND.n436 0.123142
R558 VGND.n343 VGND.n66 0.123142
R559 VGND.n438 VGND.n19 0.123127
R560 VGND.n440 VGND.n439 0.123111
R561 VGND.n443 VGND.n442 0.123081
R562 VGND.n446 VGND.n445 0.123049
R563 VGND.n402 VGND.n401 0.122488
R564 VGND.n349 VGND.n60 0.122488
R565 VGND.n435 VGND.n20 0.122394
R566 VGND.n344 VGND.n65 0.122394
R567 VGND.n287 VGND.n286 0.12129
R568 VGND.n190 VGND.n186 0.120292
R569 VGND.n194 VGND.n186 0.120292
R570 VGND.n195 VGND.n194 0.120292
R571 VGND.n196 VGND.n195 0.120292
R572 VGND.n196 VGND.n184 0.120292
R573 VGND.n184 VGND.n182 0.120292
R574 VGND.n201 VGND.n182 0.120292
R575 VGND.n202 VGND.n201 0.120292
R576 VGND.n203 VGND.n202 0.120292
R577 VGND.n203 VGND.n180 0.120292
R578 VGND.n207 VGND.n180 0.120292
R579 VGND.n208 VGND.n207 0.120292
R580 VGND.n208 VGND.n177 0.120292
R581 VGND.n212 VGND.n177 0.120292
R582 VGND.n213 VGND.n212 0.120292
R583 VGND.n214 VGND.n213 0.120292
R584 VGND.n223 VGND.n222 0.120292
R585 VGND.n223 VGND.n172 0.120292
R586 VGND.n227 VGND.n172 0.120292
R587 VGND.n228 VGND.n227 0.120292
R588 VGND.n229 VGND.n228 0.120292
R589 VGND.n229 VGND.n170 0.120292
R590 VGND.n170 VGND.n168 0.120292
R591 VGND.n234 VGND.n168 0.120292
R592 VGND.n235 VGND.n234 0.120292
R593 VGND.n236 VGND.n235 0.120292
R594 VGND.n236 VGND.n166 0.120292
R595 VGND.n166 VGND.n164 0.120292
R596 VGND.n242 VGND.n164 0.120292
R597 VGND.n243 VGND.n242 0.120292
R598 VGND.n244 VGND.n243 0.120292
R599 VGND.n244 VGND.n161 0.120292
R600 VGND.n248 VGND.n161 0.120292
R601 VGND.n312 VGND.n311 0.120292
R602 VGND.n311 VGND.n253 0.120292
R603 VGND.n307 VGND.n253 0.120292
R604 VGND.n307 VGND.n306 0.120292
R605 VGND.n306 VGND.n305 0.120292
R606 VGND.n305 VGND.n255 0.120292
R607 VGND.n301 VGND.n255 0.120292
R608 VGND.n301 VGND.n300 0.120292
R609 VGND.n300 VGND.n299 0.120292
R610 VGND.n299 VGND.n258 0.120292
R611 VGND.n259 VGND.n258 0.120292
R612 VGND.n294 VGND.n259 0.120292
R613 VGND.n294 VGND.n293 0.120292
R614 VGND.n293 VGND.n262 0.120292
R615 VGND.n289 VGND.n262 0.120292
R616 VGND.n460 VGND.n459 0.117964
R617 VGND.n375 VGND.n374 0.117514
R618 VGND.n459 VGND.n458 0.115687
R619 VGND.n458 VGND.n13 0.114144
R620 VGND.n283 VGND.n282 0.11377
R621 VGND.n454 VGND.n13 0.112073
R622 VGND.n454 VGND.n453 0.110115
R623 VGND.n374 VGND.n373 0.109841
R624 VGND.n453 VGND.n452 0.108641
R625 VGND.n452 VGND.n15 0.108047
R626 VGND.n373 VGND.n372 0.107742
R627 VGND.n339 VGND.n66 0.107432
R628 VGND.n429 VGND.n21 0.107207
R629 VGND.n448 VGND.n15 0.106987
R630 VGND.n461 VGND.n12 0.106615
R631 VGND.n448 VGND.n447 0.106444
R632 VGND.n446 VGND.n17 0.105637
R633 VGND.n447 VGND.n446 0.1051
R634 VGND.n442 VGND.n17 0.104369
R635 VGND.n457 VGND.n12 0.104071
R636 VGND.n442 VGND.n441 0.103621
R637 VGND.n123 VGND.n122 0.102649
R638 VGND.n441 VGND.n440 0.102402
R639 VGND.n457 VGND.n456 0.101564
R640 VGND.n440 VGND.n19 0.101442
R641 VGND.n436 VGND.n19 0.101268
R642 VGND.n434 VGND.n21 0.101046
R643 VGND.n346 VGND.n345 0.101046
R644 VGND.n435 VGND.n434 0.100296
R645 VGND.n345 VGND.n344 0.100296
R646 VGND.n436 VGND.n435 0.10015
R647 VGND.n344 VGND.n343 0.10015
R648 VGND.n456 VGND.n455 0.0992762
R649 VGND.n372 VGND.n371 0.0989862
R650 VGND.n222 VGND 0.0981562
R651 VGND VGND.n312 0.0981562
R652 VGND.n347 VGND.n346 0.0977333
R653 VGND.n430 VGND.n23 0.0968923
R654 VGND.n348 VGND.n347 0.0968923
R655 VGND.n125 VGND.n124 0.0967441
R656 VGND.n403 VGND.n402 0.0962186
R657 VGND.n350 VGND.n349 0.0962186
R658 VGND.n455 VGND.n14 0.0961897
R659 VGND.n402 VGND.n23 0.0958953
R660 VGND.n349 VGND.n348 0.0958953
R661 VGND.n404 VGND.n403 0.0954608
R662 VGND.n351 VGND.n350 0.0954608
R663 VGND.n108 VGND.n107 0.0953547
R664 VGND.n451 VGND.n14 0.0944655
R665 VGND.n371 VGND.n370 0.094367
R666 VGND.n370 VGND.n369 0.093816
R667 VGND.n405 VGND.n404 0.0937058
R668 VGND.n352 VGND.n351 0.0937058
R669 VGND.n462 VGND.n11 0.0936756
R670 VGND.n406 VGND.n405 0.0923613
R671 VGND.n353 VGND.n352 0.0923613
R672 VGND.n110 VGND.n109 0.0923379
R673 VGND.n109 VGND.n108 0.091697
R674 VGND.n451 VGND.n450 0.0914864
R675 VGND.n407 VGND.n406 0.091171
R676 VGND.n354 VGND.n353 0.091171
R677 VGND.n369 VGND.n368 0.0901409
R678 VGND.n409 VGND.n408 0.0898275
R679 VGND.n356 VGND.n355 0.0898275
R680 VGND.n408 VGND.n407 0.0898264
R681 VGND.n355 VGND.n354 0.0898264
R682 VGND.n343 VGND.n342 0.0897029
R683 VGND.n122 VGND.n121 0.0896537
R684 VGND.n121 VGND.n120 0.0895697
R685 VGND.n450 VGND.n449 0.0894262
R686 VGND.n113 VGND.n112 0.0883936
R687 VGND.n120 VGND.n119 0.0881488
R688 VGND.n112 VGND.n111 0.0880457
R689 VGND.n111 VGND.n110 0.0876429
R690 VGND.n116 VGND.n115 0.0874298
R691 VGND.n410 VGND.n409 0.0872535
R692 VGND.n357 VGND.n356 0.0872535
R693 VGND.n368 VGND.n367 0.0869298
R694 VGND.n449 VGND.n16 0.0869094
R695 VGND.n119 VGND.n118 0.0868534
R696 VGND.n411 VGND.n410 0.0866383
R697 VGND.n358 VGND.n357 0.0866383
R698 VGND.n114 VGND.n113 0.0862719
R699 VGND.n115 VGND.n114 0.0855718
R700 VGND.n118 VGND.n117 0.08542
R701 VGND.n367 VGND.n366 0.0853466
R702 VGND.n445 VGND.n16 0.0849371
R703 VGND.n412 VGND.n411 0.0847408
R704 VGND.n359 VGND.n358 0.0847408
R705 VGND.n117 VGND.n116 0.0846042
R706 VGND.n364 VGND.n363 0.0845436
R707 VGND.n365 VGND.n364 0.0840598
R708 VGND.n418 VGND.n417 0.0835123
R709 VGND.n366 VGND.n365 0.0835123
R710 VGND.n413 VGND.n412 0.0828145
R711 VGND.n360 VGND.n359 0.0828145
R712 VGND.n445 VGND.n444 0.0821993
R713 VGND.n416 VGND.n415 0.0819394
R714 VGND.n415 VGND.n414 0.0813683
R715 VGND.n417 VGND.n416 0.0813424
R716 VGND.n414 VGND.n413 0.0809598
R717 VGND.n444 VGND.n443 0.0805654
R718 VGND.n363 VGND.n362 0.0801429
R719 VGND.n443 VGND.n18 0.0779194
R720 VGND.n419 VGND.n418 0.0765448
R721 VGND.n439 VGND.n18 0.0763064
R722 VGND.n189 VGND 0.0758148
R723 VGND.n125 VGND.n79 0.0740294
R724 VGND.n439 VGND.n438 0.0737484
R725 VGND.n438 VGND.n437 0.0717025
R726 VGND.n437 VGND.n20 0.0696824
R727 VGND.n66 VGND.n65 0.0696824
R728 VGND.n361 VGND.n360 0.0694343
R729 VGND.n433 VGND.n20 0.0672702
R730 VGND.n65 VGND.n64 0.0672702
R731 VGND.n433 VGND.n432 0.0664938
R732 VGND.n64 VGND.n63 0.0664938
R733 VGND.n432 VGND.n431 0.0637716
R734 VGND.n63 VGND.n62 0.0637716
R735 VGND.n431 VGND.n22 0.0618497
R736 VGND.n62 VGND.n61 0.0618497
R737 VGND.n419 VGND.n384 0.0612585
R738 VGND.n214 VGND 0.0603958
R739 VGND.n217 VGND 0.0603958
R740 VGND.n218 VGND 0.0603958
R741 VGND.n221 VGND 0.0603958
R742 VGND VGND.n248 0.0603958
R743 VGND.n249 VGND 0.0603958
R744 VGND.n250 VGND 0.0603958
R745 VGND.n313 VGND 0.0603958
R746 VGND.n401 VGND.n22 0.0599512
R747 VGND.n61 VGND.n60 0.0599512
R748 VGND.n401 VGND.n400 0.0577289
R749 VGND.n60 VGND.n59 0.0577289
R750 VGND.n48 VGND 0.05675
R751 VGND.n337 VGND 0.05675
R752 VGND.n146 VGND 0.05675
R753 VGND.n428 VGND 0.05675
R754 VGND.n10 VGND 0.05675
R755 VGND.n467 VGND 0.05675
R756 VGND.n326 VGND 0.05675
R757 VGND.n341 VGND 0.05675
R758 VGND.n319 VGND 0.05675
R759 VGND.n420 VGND 0.05675
R760 VGND.n400 VGND.n399 0.0562229
R761 VGND.n59 VGND.n58 0.0562229
R762 VGND.n399 VGND.n398 0.0543922
R763 VGND.n58 VGND.n57 0.0543922
R764 VGND.n460 VGND.n11 0.0535576
R765 VGND.n398 VGND.n397 0.0525833
R766 VGND.n57 VGND.n56 0.0525833
R767 VGND.n80 VGND.n79 0.0506497
R768 VGND.n397 VGND.n396 0.0503512
R769 VGND.n56 VGND.n55 0.0503512
R770 VGND.n385 VGND.n384 0.0500244
R771 VGND.n81 VGND.n80 0.0496071
R772 VGND.n477 VGND.n1 0.0495625
R773 VGND.n396 VGND.n395 0.0490294
R774 VGND.n55 VGND.n54 0.0490294
R775 VGND.n342 VGND.n339 0.0489751
R776 VGND.n82 VGND.n81 0.047375
R777 VGND.n395 VGND.n394 0.0468235
R778 VGND.n54 VGND.n53 0.0468235
R779 VGND.n83 VGND.n82 0.0460882
R780 VGND.n394 VGND.n393 0.0458216
R781 VGND.n53 VGND.n52 0.0458216
R782 VGND.n84 VGND.n83 0.0438824
R783 VGND.n393 VGND.n392 0.0433779
R784 VGND.n52 VGND.n51 0.0433779
R785 VGND.n126 VGND.n125 0.0427535
R786 VGND.n85 VGND.n84 0.0421667
R787 VGND.n392 VGND.n391 0.0419244
R788 VGND.n51 VGND.n50 0.0419244
R789 VGND.n86 VGND.n85 0.0404709
R790 VGND.n391 VGND.n390 0.0402399
R791 VGND.n50 VGND.n49 0.0402399
R792 VGND.n87 VGND.n86 0.0382907
R793 VGND.n390 VGND.n389 0.0378563
R794 VGND.n49 VGND.n47 0.0378563
R795 VGND.n88 VGND.n87 0.0373497
R796 VGND.n389 VGND.n388 0.0371379
R797 VGND.n47 VGND.n46 0.0371379
R798 VGND.n89 VGND.n88 0.0349828
R799 VGND.n388 VGND.n387 0.0347857
R800 VGND.n46 VGND.n45 0.0347857
R801 VGND VGND.n217 0.0343542
R802 VGND.n218 VGND 0.0343542
R803 VGND VGND.n249 0.0343542
R804 VGND VGND.n250 0.0343542
R805 VGND.n90 VGND.n89 0.033546
R806 VGND.n387 VGND.n386 0.0331705
R807 VGND.n45 VGND.n44 0.0331705
R808 VGND.n91 VGND.n90 0.0319286
R809 VGND.n386 VGND.n385 0.03175
R810 VGND.n44 VGND.n43 0.03175
R811 VGND.n126 VGND.n2 0.0315536
R812 VGND.n430 VGND.n429 0.0311748
R813 VGND.n92 VGND.n91 0.0303295
R814 VGND.n43 VGND.n42 0.030161
R815 VGND.n478 VGND.n0 0.0288333
R816 VGND.n479 VGND.n478 0.0288333
R817 VGND.n93 VGND.n92 0.0281989
R818 VGND.n42 VGND.n41 0.0280424
R819 VGND.n94 VGND.n93 0.0266299
R820 VGND.n41 VGND.n40 0.0266299
R821 VGND.n95 VGND.n94 0.0252175
R822 VGND.n40 VGND.n39 0.0250787
R823 VGND.n105 VGND.n95 0.0238051
R824 VGND.n39 VGND.n38 0.0235447
R825 VGND VGND.n221 0.0226354
R826 VGND.n313 VGND 0.0226354
R827 VGND.n38 VGND.n37 0.0222697
R828 VGND.n37 VGND.n36 0.0200531
R829 VGND.n36 VGND.n35 0.0185556
R830 VGND.n35 VGND.n34 0.0172598
R831 VGND.n284 VGND.n283 0.01695
R832 VGND.n34 VGND.n33 0.0157778
R833 VGND.n362 VGND.n361 0.0153586
R834 VGND.n33 VGND.n32 0.0136944
R835 VGND.n106 VGND.n105 0.0123255
R836 VGND.n32 VGND.n31 0.0122403
R837 VGND.n31 VGND.n30 0.0109167
R838 VGND.n287 VGND.n272 0.00943
R839 VGND.n30 VGND.n29 0.00878729
R840 VGND.n383 VGND.n382 0.00778193
R841 VGND.n382 VGND.n29 0.00740608
R842 VAPWR.n52 VAPWR.t13 738.799
R843 VAPWR.n50 VAPWR.t21 738.799
R844 VAPWR.n23 VAPWR.t19 738.799
R845 VAPWR.n16 VAPWR.t27 738.799
R846 VAPWR.n15 VAPWR.t5 738.799
R847 VAPWR.n100 VAPWR.t7 738.799
R848 VAPWR.n17 VAPWR.t11 738.799
R849 VAPWR.n18 VAPWR.t15 738.799
R850 VAPWR.n21 VAPWR.t9 738.799
R851 VAPWR.n25 VAPWR.t17 738.799
R852 VAPWR.n48 VAPWR.t41 738.799
R853 VAPWR.n0 VAPWR.t29 738.799
R854 VAPWR.n84 VAPWR.t35 738.799
R855 VAPWR.n13 VAPWR.t3 738.799
R856 VAPWR.n5 VAPWR.t31 738.799
R857 VAPWR.n3 VAPWR.t33 738.799
R858 VAPWR.n97 VAPWR.t37 738.799
R859 VAPWR.n7 VAPWR.t39 738.799
R860 VAPWR.n9 VAPWR.t1 738.799
R861 VAPWR.n11 VAPWR.t23 738.799
R862 VAPWR.n89 VAPWR.t25 738.799
R863 VAPWR.n0 VAPWR.t28 707.519
R864 VAPWR.n52 VAPWR.t12 707.519
R865 VAPWR.n50 VAPWR.t20 707.519
R866 VAPWR.n23 VAPWR.t18 707.519
R867 VAPWR.n16 VAPWR.t26 707.519
R868 VAPWR.n84 VAPWR.t34 707.519
R869 VAPWR.n15 VAPWR.t4 707.519
R870 VAPWR.n13 VAPWR.t2 707.519
R871 VAPWR.n5 VAPWR.t30 707.519
R872 VAPWR.n3 VAPWR.t32 707.519
R873 VAPWR.n97 VAPWR.t36 707.519
R874 VAPWR.n100 VAPWR.t6 707.519
R875 VAPWR.n7 VAPWR.t38 707.519
R876 VAPWR.n9 VAPWR.t0 707.519
R877 VAPWR.n11 VAPWR.t22 707.519
R878 VAPWR.n89 VAPWR.t24 707.519
R879 VAPWR.n17 VAPWR.t10 707.519
R880 VAPWR.n18 VAPWR.t14 707.519
R881 VAPWR.n21 VAPWR.t8 707.519
R882 VAPWR.n25 VAPWR.t16 707.519
R883 VAPWR.n48 VAPWR.t40 707.519
R884 VAPWR.n1 VAPWR.n0 13.3797
R885 VAPWR.n85 VAPWR.n84 13.3797
R886 VAPWR.n14 VAPWR.n13 13.3797
R887 VAPWR.n6 VAPWR.n5 13.3797
R888 VAPWR.n4 VAPWR.n3 13.3797
R889 VAPWR.n98 VAPWR.n97 13.3797
R890 VAPWR.n8 VAPWR.n7 13.3797
R891 VAPWR.n10 VAPWR.n9 13.3797
R892 VAPWR.n12 VAPWR.n11 13.3797
R893 VAPWR.n90 VAPWR.n89 13.3797
R894 VAPWR VAPWR.n52 13.3223
R895 VAPWR.n51 VAPWR.n50 13.3223
R896 VAPWR.n24 VAPWR.n23 13.3223
R897 VAPWR VAPWR.n16 13.3223
R898 VAPWR VAPWR.n15 13.3223
R899 VAPWR VAPWR.n100 13.3223
R900 VAPWR VAPWR.n17 13.3223
R901 VAPWR.n19 VAPWR.n18 13.3223
R902 VAPWR.n22 VAPWR.n21 13.3223
R903 VAPWR.n26 VAPWR.n25 13.3223
R904 VAPWR.n49 VAPWR.n48 13.3223
R905 VAPWR.n83 VAPWR.n82 13.3027
R906 VAPWR.n53 VAPWR 12.2181
R907 VAPWR.n83 VAPWR 9.41984
R908 VAPWR.n2 VAPWR.n1 8.84871
R909 VAPWR.n20 VAPWR 8.23756
R910 VAPWR.n87 VAPWR 7.89226
R911 VAPWR.n99 VAPWR.n98 7.80052
R912 VAPWR.n92 VAPWR.n91 7.55311
R913 VAPWR.n96 VAPWR.n4 7.50807
R914 VAPWR.n86 VAPWR.n85 7.20658
R915 VAPWR.n101 VAPWR 7.08652
R916 VAPWR.n95 VAPWR.n6 6.80411
R917 VAPWR.n91 VAPWR.n88 6.76495
R918 VAPWR.n54 VAPWR.n51 6.56755
R919 VAPWR.n81 VAPWR.n22 6.51187
R920 VAPWR.n88 VAPWR.n14 6.43822
R921 VAPWR.n99 VAPWR.n96 6.22803
R922 VAPWR.n94 VAPWR.n8 6.22106
R923 VAPWR.n80 VAPWR.n24 6.09916
R924 VAPWR.n91 VAPWR.n90 6.0818
R925 VAPWR.n93 VAPWR.n10 6.01232
R926 VAPWR.n92 VAPWR.n12 5.93615
R927 VAPWR.n56 VAPWR.n49 5.89109
R928 VAPWR.n27 VAPWR.n26 5.80982
R929 VAPWR.n20 VAPWR.n19 4.80965
R930 VAPWR.n95 VAPWR.n94 4.15423
R931 VAPWR.n53 VAPWR.n2 3.74435
R932 VAPWR.n103 VAPWR 3.46747
R933 VAPWR.n104 VAPWR 3.41928
R934 VAPWR.n54 VAPWR.n53 3.13707
R935 VAPWR.n96 VAPWR.n95 2.87981
R936 VAPWR.n82 VAPWR.n20 2.79302
R937 VAPWR.n103 VAPWR.n102 1.13771
R938 VAPWR.n101 VAPWR.n99 1.13693
R939 VAPWR.n93 VAPWR.n92 0.937335
R940 VAPWR.n87 VAPWR.n86 0.929914
R941 VAPWR.n81 VAPWR.n80 0.915244
R942 VAPWR.n86 VAPWR.n83 0.904418
R943 VAPWR.n55 VAPWR.n54 0.893623
R944 VAPWR.n94 VAPWR.n93 0.872816
R945 VAPWR.n102 VAPWR.n2 0.848313
R946 VAPWR.n88 VAPWR.n87 0.756987
R947 VAPWR.n80 VAPWR.n79 0.51791
R948 VAPWR.n79 VAPWR.n27 0.319334
R949 VAPWR.n82 VAPWR.n81 0.302419
R950 VAPWR VAPWR.n104 0.190997
R951 VAPWR.n58 VAPWR.n57 0.153341
R952 VAPWR.n55 VAPWR.n47 0.138117
R953 VAPWR.n76 VAPWR.n28 0.136106
R954 VAPWR.n78 VAPWR.n77 0.136042
R955 VAPWR.n73 VAPWR.n31 0.135531
R956 VAPWR.n74 VAPWR.n30 0.135469
R957 VAPWR.n75 VAPWR.n29 0.135409
R958 VAPWR.n58 VAPWR.n46 0.135115
R959 VAPWR.n59 VAPWR.n45 0.135049
R960 VAPWR.n70 VAPWR.n34 0.134934
R961 VAPWR.n60 VAPWR.n44 0.134918
R962 VAPWR.n61 VAPWR.n43 0.134854
R963 VAPWR.n72 VAPWR.n32 0.134817
R964 VAPWR.n62 VAPWR.n42 0.134728
R965 VAPWR.n64 VAPWR.n40 0.134606
R966 VAPWR.n65 VAPWR.n39 0.134487
R967 VAPWR.n67 VAPWR.n37 0.134371
R968 VAPWR.n69 VAPWR.n35 0.134203
R969 VAPWR.n63 VAPWR.n41 0.133778
R970 VAPWR.n66 VAPWR.n38 0.133565
R971 VAPWR.n68 VAPWR.n36 0.133462
R972 VAPWR.n71 VAPWR.n33 0.133264
R973 VAPWR.n77 VAPWR.n76 0.122659
R974 VAPWR.n76 VAPWR.n75 0.122197
R975 VAPWR.n60 VAPWR.n59 0.117149
R976 VAPWR.n59 VAPWR.n58 0.117099
R977 VAPWR.n75 VAPWR.n74 0.116731
R978 VAPWR.n61 VAPWR.n60 0.114696
R979 VAPWR.n73 VAPWR.n72 0.1146
R980 VAPWR.n74 VAPWR.n73 0.114178
R981 VAPWR.n62 VAPWR.n61 0.113375
R982 VAPWR.n72 VAPWR.n71 0.113293
R983 VAPWR.n63 VAPWR.n62 0.111589
R984 VAPWR.n65 VAPWR.n64 0.110724
R985 VAPWR.n64 VAPWR.n63 0.110707
R986 VAPWR.n69 VAPWR.n68 0.110107
R987 VAPWR.n70 VAPWR.n69 0.109771
R988 VAPWR.n67 VAPWR.n66 0.109608
R989 VAPWR.n68 VAPWR.n67 0.109359
R990 VAPWR.n66 VAPWR.n65 0.109137
R991 VAPWR.n71 VAPWR.n70 0.10735
R992 VAPWR.n57 VAPWR.n47 0.0846195
R993 VAPWR.n47 VAPWR.n46 0.0809196
R994 VAPWR.n46 VAPWR.n45 0.078625
R995 VAPWR.n45 VAPWR.n44 0.0749863
R996 VAPWR.n56 VAPWR.n55 0.0739204
R997 VAPWR.n44 VAPWR.n43 0.0719286
R998 VAPWR.n43 VAPWR.n42 0.068453
R999 VAPWR.n42 VAPWR.n41 0.0658974
R1000 VAPWR.n41 VAPWR.n40 0.0642417
R1001 VAPWR.n40 VAPWR.n39 0.0601405
R1002 VAPWR.n57 VAPWR.n56 0.057945
R1003 VAPWR.n1 VAPWR 0.057877
R1004 VAPWR.n85 VAPWR 0.057877
R1005 VAPWR.n14 VAPWR 0.057877
R1006 VAPWR.n6 VAPWR 0.057877
R1007 VAPWR.n4 VAPWR 0.057877
R1008 VAPWR.n98 VAPWR 0.057877
R1009 VAPWR.n8 VAPWR 0.057877
R1010 VAPWR.n10 VAPWR 0.057877
R1011 VAPWR.n12 VAPWR 0.057877
R1012 VAPWR.n90 VAPWR 0.057877
R1013 VAPWR.n39 VAPWR.n38 0.0577581
R1014 VAPWR.n38 VAPWR.n37 0.0553387
R1015 VAPWR.n37 VAPWR.n36 0.0530478
R1016 VAPWR.n36 VAPWR.n35 0.0503418
R1017 VAPWR.n51 VAPWR 0.0496071
R1018 VAPWR.n24 VAPWR 0.0496071
R1019 VAPWR.n19 VAPWR 0.0496071
R1020 VAPWR.n22 VAPWR 0.0496071
R1021 VAPWR.n26 VAPWR 0.0496071
R1022 VAPWR.n49 VAPWR 0.0496071
R1023 VAPWR.n35 VAPWR.n34 0.0468836
R1024 VAPWR.n34 VAPWR.n33 0.0455311
R1025 VAPWR.n33 VAPWR.n32 0.0424255
R1026 VAPWR.n79 VAPWR.n78 0.042321
R1027 VAPWR.n32 VAPWR.n31 0.0398519
R1028 VAPWR.n31 VAPWR.n30 0.0380767
R1029 VAPWR.n30 VAPWR.n29 0.035561
R1030 VAPWR.n29 VAPWR.n28 0.0323182
R1031 VAPWR.n78 VAPWR.n28 0.0306205
R1032 VAPWR.n102 VAPWR.n101 0.0273117
R1033 VAPWR.n77 VAPWR.n27 0.0155602
R1034 VAPWR.n104 VAPWR.n103 0.00193165
R1035 uo_out[2].n2 uo_out[2].t1 313.104
R1036 uo_out[2].n0 uo_out[2].t2 294.557
R1037 uo_out[2].t0 uo_out[2].n2 265.769
R1038 uo_out[2] uo_out[2].t0 262.318
R1039 uo_out[2].n0 uo_out[2].t3 211.01
R1040 uo_out[2].n1 uo_out[2].n0 152
R1041 uo_out[2].n5 uo_out[2] 16.2155
R1042 uo_out[2].n4 uo_out[2].n1 11.6311
R1043 uo_out[2].n4 uo_out[2].n3 9.3005
R1044 uo_out[2].n3 uo_out[2] 7.17626
R1045 uo_out[2].n3 uo_out[2].n2 4.84898
R1046 uo_out[2].n5 uo_out[2].n4 4.51042
R1047 uo_out[2].n1 uo_out[2] 1.37896
R1048 uo_out[2] uo_out[2].n5 0.0730806
R1049 VDPWR.n1 VDPWR.t51 738.801
R1050 VDPWR.n1 VDPWR.t50 707.519
R1051 VDPWR.n84 VDPWR.t37 667.734
R1052 VDPWR.n52 VDPWR.t71 667.734
R1053 VDPWR.n124 VDPWR.t19 667.734
R1054 VDPWR.n99 VDPWR.t65 666.677
R1055 VDPWR.n38 VDPWR.t55 666.677
R1056 VDPWR.n4 VDPWR.t57 666.677
R1057 VDPWR.t46 VDPWR.t18 624.456
R1058 VDPWR.t70 VDPWR.t30 624.456
R1059 VDPWR.t36 VDPWR.t52 624.456
R1060 VDPWR.n102 VDPWR.n101 604.394
R1061 VDPWR.n33 VDPWR.n32 604.394
R1062 VDPWR.n142 VDPWR.n141 604.394
R1063 VDPWR.t56 VDPWR.t10 556.386
R1064 VDPWR.t16 VDPWR.t14 556.386
R1065 VDPWR.t60 VDPWR.t54 556.386
R1066 VDPWR.t68 VDPWR.t66 556.386
R1067 VDPWR.t24 VDPWR.t64 556.386
R1068 VDPWR.t34 VDPWR.t38 556.386
R1069 VDPWR.n17 VDPWR.t32 414.33
R1070 VDPWR.t44 VDPWR.n108 414.33
R1071 VDPWR.t42 VDPWR.t6 390.654
R1072 VDPWR.t0 VDPWR.t20 390.654
R1073 VDPWR.t28 VDPWR.t2 390.654
R1074 VDPWR.t18 VDPWR.t49 337.384
R1075 VDPWR.t5 VDPWR.t70 337.384
R1076 VDPWR.t8 VDPWR.t36 337.384
R1077 VDPWR.n82 VDPWR.n72 333.348
R1078 VDPWR.n54 VDPWR.n24 333.348
R1079 VDPWR.n122 VDPWR.n12 333.348
R1080 VDPWR.n68 VDPWR.n67 320.976
R1081 VDPWR.n45 VDPWR.n28 320.976
R1082 VDPWR.n9 VDPWR.n8 320.976
R1083 VDPWR.t6 VDPWR.t12 304.829
R1084 VDPWR.t62 VDPWR.t0 304.829
R1085 VDPWR.t22 VDPWR.t28 304.829
R1086 VDPWR.t32 VDPWR.t16 287.072
R1087 VDPWR.t66 VDPWR.t44 287.072
R1088 VDPWR.t38 VDPWR.t40 287.072
R1089 VDPWR.t12 VDPWR.t48 281.154
R1090 VDPWR.t13 VDPWR.t42 281.154
R1091 VDPWR.t4 VDPWR.t62 281.154
R1092 VDPWR.t20 VDPWR.t63 281.154
R1093 VDPWR.t9 VDPWR.t22 281.154
R1094 VDPWR.t2 VDPWR.t23 281.154
R1095 VDPWR.n109 VDPWR.n17 272.274
R1096 VDPWR.n109 VDPWR 272.274
R1097 VDPWR.n108 VDPWR.n107 272.274
R1098 VDPWR.n107 VDPWR 272.274
R1099 VDPWR.t48 VDPWR.t56 251.559
R1100 VDPWR.t54 VDPWR.t4 251.559
R1101 VDPWR.t64 VDPWR.t9 251.559
R1102 VDPWR.t10 VDPWR.t72 248.599
R1103 VDPWR.t49 VDPWR.t13 248.599
R1104 VDPWR.t14 VDPWR.t46 248.599
R1105 VDPWR.t26 VDPWR.t60 248.599
R1106 VDPWR.t63 VDPWR.t5 248.599
R1107 VDPWR.t30 VDPWR.t68 248.599
R1108 VDPWR.t58 VDPWR.t24 248.599
R1109 VDPWR.t23 VDPWR.t8 248.599
R1110 VDPWR.t52 VDPWR.t34 248.599
R1111 VDPWR.n76 VDPWR.n75 240.522
R1112 VDPWR.n60 VDPWR.n21 240.522
R1113 VDPWR.n116 VDPWR.n115 240.522
R1114 VDPWR.n107 VDPWR.n106 213.119
R1115 VDPWR.n108 VDPWR.n18 213.119
R1116 VDPWR.n110 VDPWR.n109 213.119
R1117 VDPWR.n17 VDPWR.n15 213.119
R1118 VDPWR.n67 VDPWR.t29 113.98
R1119 VDPWR.n28 VDPWR.t1 113.98
R1120 VDPWR.n8 VDPWR.t7 113.98
R1121 VDPWR.t72 VDPWR 91.745
R1122 VDPWR VDPWR.t26 91.745
R1123 VDPWR VDPWR.t58 91.745
R1124 VDPWR.n75 VDPWR.t39 61.9872
R1125 VDPWR.n21 VDPWR.t67 61.9872
R1126 VDPWR.n115 VDPWR.t17 61.9872
R1127 VDPWR.n101 VDPWR.t59 41.5552
R1128 VDPWR.n101 VDPWR.t25 41.5552
R1129 VDPWR.n32 VDPWR.t27 41.5552
R1130 VDPWR.n32 VDPWR.t61 41.5552
R1131 VDPWR.n141 VDPWR.t73 41.5552
R1132 VDPWR.n141 VDPWR.t11 41.5552
R1133 VDPWR.n67 VDPWR.t3 35.4605
R1134 VDPWR.n28 VDPWR.t21 35.4605
R1135 VDPWR.n8 VDPWR.t43 35.4605
R1136 VDPWR.n81 VDPWR.n73 34.6358
R1137 VDPWR.n77 VDPWR.n73 34.6358
R1138 VDPWR.n95 VDPWR.n65 34.6358
R1139 VDPWR.n95 VDPWR.n94 34.6358
R1140 VDPWR.n94 VDPWR.n93 34.6358
R1141 VDPWR.n90 VDPWR.n89 34.6358
R1142 VDPWR.n89 VDPWR.n88 34.6358
R1143 VDPWR.n88 VDPWR.n70 34.6358
R1144 VDPWR.n55 VDPWR.n22 34.6358
R1145 VDPWR.n59 VDPWR.n22 34.6358
R1146 VDPWR.n40 VDPWR.n39 34.6358
R1147 VDPWR.n40 VDPWR.n29 34.6358
R1148 VDPWR.n44 VDPWR.n29 34.6358
R1149 VDPWR.n47 VDPWR.n46 34.6358
R1150 VDPWR.n47 VDPWR.n26 34.6358
R1151 VDPWR.n51 VDPWR.n26 34.6358
R1152 VDPWR.n121 VDPWR.n13 34.6358
R1153 VDPWR.n117 VDPWR.n13 34.6358
R1154 VDPWR.n136 VDPWR.n135 34.6358
R1155 VDPWR.n135 VDPWR.n134 34.6358
R1156 VDPWR.n134 VDPWR.n6 34.6358
R1157 VDPWR.n130 VDPWR.n129 34.6358
R1158 VDPWR.n129 VDPWR.n128 34.6358
R1159 VDPWR.n128 VDPWR.n10 34.6358
R1160 VDPWR.n83 VDPWR.n82 32.0005
R1161 VDPWR.n54 VDPWR.n53 32.0005
R1162 VDPWR.n123 VDPWR.n122 32.0005
R1163 VDPWR.n143 VDPWR.n142 30.7593
R1164 VDPWR.n84 VDPWR.n83 30.4946
R1165 VDPWR.n53 VDPWR.n52 30.4946
R1166 VDPWR.n124 VDPWR.n123 30.4946
R1167 VDPWR.n75 VDPWR.t41 30.1692
R1168 VDPWR.n21 VDPWR.t45 30.1692
R1169 VDPWR.n115 VDPWR.t33 30.1692
R1170 VDPWR.n99 VDPWR.n65 27.4829
R1171 VDPWR.n61 VDPWR.n60 27.4829
R1172 VDPWR.n39 VDPWR.n38 27.4829
R1173 VDPWR.n116 VDPWR.n114 27.4829
R1174 VDPWR.n136 VDPWR.n4 27.4829
R1175 VDPWR.n72 VDPWR.t53 26.5955
R1176 VDPWR.n72 VDPWR.t35 26.5955
R1177 VDPWR.n24 VDPWR.t31 26.5955
R1178 VDPWR.n24 VDPWR.t69 26.5955
R1179 VDPWR.n12 VDPWR.t47 26.5955
R1180 VDPWR.n12 VDPWR.t15 26.5955
R1181 VDPWR.n77 VDPWR.n76 25.6005
R1182 VDPWR.n60 VDPWR.n59 25.6005
R1183 VDPWR.n117 VDPWR.n116 25.6005
R1184 VDPWR.n106 VDPWR.n19 23.7181
R1185 VDPWR.n61 VDPWR.n18 23.7181
R1186 VDPWR.n110 VDPWR.n16 23.7181
R1187 VDPWR.n114 VDPWR.n15 23.7181
R1188 VDPWR.n102 VDPWR.n100 22.9652
R1189 VDPWR.n37 VDPWR.n33 22.9652
R1190 VDPWR.n142 VDPWR.n140 22.9652
R1191 VDPWR.n100 VDPWR.n99 21.8358
R1192 VDPWR.n38 VDPWR.n37 21.8358
R1193 VDPWR.n140 VDPWR.n4 21.8358
R1194 VDPWR.n102 VDPWR.n19 21.4593
R1195 VDPWR.n33 VDPWR.n16 21.4593
R1196 VDPWR.n93 VDPWR.n68 18.4476
R1197 VDPWR.n45 VDPWR.n44 18.4476
R1198 VDPWR.n9 VDPWR.n6 18.4476
R1199 VDPWR.n90 VDPWR.n68 16.1887
R1200 VDPWR.n46 VDPWR.n45 16.1887
R1201 VDPWR.n130 VDPWR.n9 16.1887
R1202 VDPWR.n84 VDPWR.n70 15.0593
R1203 VDPWR.n52 VDPWR.n51 15.0593
R1204 VDPWR.n124 VDPWR.n10 15.0593
R1205 VDPWR.n2 VDPWR.n1 13.3223
R1206 VDPWR.n106 VDPWR.n18 12.8005
R1207 VDPWR.n110 VDPWR.n15 12.8005
R1208 VDPWR.n3 VDPWR 10.4749
R1209 VDPWR.n143 VDPWR.n3 9.61724
R1210 VDPWR.n142 VDPWR.n0 9.3005
R1211 VDPWR.n140 VDPWR.n139 9.3005
R1212 VDPWR.n138 VDPWR.n4 9.3005
R1213 VDPWR.n137 VDPWR.n136 9.3005
R1214 VDPWR.n135 VDPWR.n5 9.3005
R1215 VDPWR.n134 VDPWR.n133 9.3005
R1216 VDPWR.n132 VDPWR.n6 9.3005
R1217 VDPWR.n131 VDPWR.n130 9.3005
R1218 VDPWR.n129 VDPWR.n7 9.3005
R1219 VDPWR.n128 VDPWR.n127 9.3005
R1220 VDPWR.n126 VDPWR.n10 9.3005
R1221 VDPWR.n125 VDPWR.n124 9.3005
R1222 VDPWR.n123 VDPWR.n11 9.3005
R1223 VDPWR.n121 VDPWR.n120 9.3005
R1224 VDPWR.n119 VDPWR.n13 9.3005
R1225 VDPWR.n118 VDPWR.n117 9.3005
R1226 VDPWR.n116 VDPWR.n14 9.3005
R1227 VDPWR.n114 VDPWR.n113 9.3005
R1228 VDPWR.n112 VDPWR.n15 9.3005
R1229 VDPWR.n111 VDPWR.n110 9.3005
R1230 VDPWR.n34 VDPWR.n16 9.3005
R1231 VDPWR.n35 VDPWR.n33 9.3005
R1232 VDPWR.n37 VDPWR.n36 9.3005
R1233 VDPWR.n38 VDPWR.n31 9.3005
R1234 VDPWR.n39 VDPWR.n30 9.3005
R1235 VDPWR.n41 VDPWR.n40 9.3005
R1236 VDPWR.n42 VDPWR.n29 9.3005
R1237 VDPWR.n44 VDPWR.n43 9.3005
R1238 VDPWR.n46 VDPWR.n27 9.3005
R1239 VDPWR.n48 VDPWR.n47 9.3005
R1240 VDPWR.n49 VDPWR.n26 9.3005
R1241 VDPWR.n51 VDPWR.n50 9.3005
R1242 VDPWR.n52 VDPWR.n25 9.3005
R1243 VDPWR.n53 VDPWR.n23 9.3005
R1244 VDPWR.n56 VDPWR.n55 9.3005
R1245 VDPWR.n57 VDPWR.n22 9.3005
R1246 VDPWR.n59 VDPWR.n58 9.3005
R1247 VDPWR.n60 VDPWR.n20 9.3005
R1248 VDPWR.n62 VDPWR.n61 9.3005
R1249 VDPWR.n63 VDPWR.n18 9.3005
R1250 VDPWR.n106 VDPWR.n105 9.3005
R1251 VDPWR.n104 VDPWR.n19 9.3005
R1252 VDPWR.n103 VDPWR.n102 9.3005
R1253 VDPWR.n100 VDPWR.n64 9.3005
R1254 VDPWR.n99 VDPWR.n98 9.3005
R1255 VDPWR.n97 VDPWR.n65 9.3005
R1256 VDPWR.n96 VDPWR.n95 9.3005
R1257 VDPWR.n94 VDPWR.n66 9.3005
R1258 VDPWR.n93 VDPWR.n92 9.3005
R1259 VDPWR.n91 VDPWR.n90 9.3005
R1260 VDPWR.n89 VDPWR.n69 9.3005
R1261 VDPWR.n88 VDPWR.n87 9.3005
R1262 VDPWR.n86 VDPWR.n70 9.3005
R1263 VDPWR.n85 VDPWR.n84 9.3005
R1264 VDPWR.n83 VDPWR.n71 9.3005
R1265 VDPWR.n81 VDPWR.n80 9.3005
R1266 VDPWR.n79 VDPWR.n73 9.3005
R1267 VDPWR.n78 VDPWR.n77 9.3005
R1268 VDPWR.n3 VDPWR.n2 8.39487
R1269 VDPWR.n76 VDPWR.n74 7.4049
R1270 VDPWR.n82 VDPWR.n81 2.63579
R1271 VDPWR.n55 VDPWR.n54 2.63579
R1272 VDPWR.n122 VDPWR.n121 2.63579
R1273 VDPWR.n74 VDPWR 0.156264
R1274 VDPWR.n78 VDPWR.n74 0.144904
R1275 VDPWR.n139 VDPWR.n0 0.120292
R1276 VDPWR.n139 VDPWR.n138 0.120292
R1277 VDPWR.n138 VDPWR.n137 0.120292
R1278 VDPWR.n137 VDPWR.n5 0.120292
R1279 VDPWR.n133 VDPWR.n5 0.120292
R1280 VDPWR.n133 VDPWR.n132 0.120292
R1281 VDPWR.n132 VDPWR.n131 0.120292
R1282 VDPWR.n131 VDPWR.n7 0.120292
R1283 VDPWR.n127 VDPWR.n7 0.120292
R1284 VDPWR.n127 VDPWR.n126 0.120292
R1285 VDPWR.n126 VDPWR.n125 0.120292
R1286 VDPWR.n125 VDPWR.n11 0.120292
R1287 VDPWR.n120 VDPWR.n11 0.120292
R1288 VDPWR.n120 VDPWR.n119 0.120292
R1289 VDPWR.n119 VDPWR.n118 0.120292
R1290 VDPWR.n118 VDPWR.n14 0.120292
R1291 VDPWR.n113 VDPWR.n14 0.120292
R1292 VDPWR.n36 VDPWR.n35 0.120292
R1293 VDPWR.n36 VDPWR.n31 0.120292
R1294 VDPWR.n31 VDPWR.n30 0.120292
R1295 VDPWR.n41 VDPWR.n30 0.120292
R1296 VDPWR.n42 VDPWR.n41 0.120292
R1297 VDPWR.n43 VDPWR.n42 0.120292
R1298 VDPWR.n43 VDPWR.n27 0.120292
R1299 VDPWR.n48 VDPWR.n27 0.120292
R1300 VDPWR.n49 VDPWR.n48 0.120292
R1301 VDPWR.n50 VDPWR.n49 0.120292
R1302 VDPWR.n50 VDPWR.n25 0.120292
R1303 VDPWR.n25 VDPWR.n23 0.120292
R1304 VDPWR.n56 VDPWR.n23 0.120292
R1305 VDPWR.n57 VDPWR.n56 0.120292
R1306 VDPWR.n58 VDPWR.n57 0.120292
R1307 VDPWR.n58 VDPWR.n20 0.120292
R1308 VDPWR.n62 VDPWR.n20 0.120292
R1309 VDPWR.n103 VDPWR.n64 0.120292
R1310 VDPWR.n98 VDPWR.n64 0.120292
R1311 VDPWR.n98 VDPWR.n97 0.120292
R1312 VDPWR.n97 VDPWR.n96 0.120292
R1313 VDPWR.n96 VDPWR.n66 0.120292
R1314 VDPWR.n92 VDPWR.n66 0.120292
R1315 VDPWR.n92 VDPWR.n91 0.120292
R1316 VDPWR.n91 VDPWR.n69 0.120292
R1317 VDPWR.n87 VDPWR.n69 0.120292
R1318 VDPWR.n87 VDPWR.n86 0.120292
R1319 VDPWR.n86 VDPWR.n85 0.120292
R1320 VDPWR.n85 VDPWR.n71 0.120292
R1321 VDPWR.n80 VDPWR.n71 0.120292
R1322 VDPWR.n80 VDPWR.n79 0.120292
R1323 VDPWR.n79 VDPWR.n78 0.120292
R1324 VDPWR VDPWR.n0 0.0981562
R1325 VDPWR.n35 VDPWR 0.0981562
R1326 VDPWR VDPWR.n103 0.0981562
R1327 VDPWR.n113 VDPWR 0.0603958
R1328 VDPWR VDPWR.n112 0.0603958
R1329 VDPWR VDPWR.n111 0.0603958
R1330 VDPWR.n34 VDPWR 0.0603958
R1331 VDPWR VDPWR.n62 0.0603958
R1332 VDPWR.n63 VDPWR 0.0603958
R1333 VDPWR.n105 VDPWR 0.0603958
R1334 VDPWR VDPWR.n104 0.0603958
R1335 VDPWR.n2 VDPWR 0.0496071
R1336 VDPWR.n112 VDPWR 0.0382604
R1337 VDPWR.n111 VDPWR 0.0382604
R1338 VDPWR VDPWR.n63 0.0382604
R1339 VDPWR.n105 VDPWR 0.0382604
R1340 VDPWR VDPWR.n34 0.0226354
R1341 VDPWR.n104 VDPWR 0.0226354
R1342 VDPWR VDPWR.n143 0.0224072
R1343 uo_out[1].n2 uo_out[1].t0 313.104
R1344 uo_out[1].n0 uo_out[1].t2 294.557
R1345 uo_out[1].t1 uo_out[1].n2 265.769
R1346 uo_out[1] uo_out[1].t1 262.318
R1347 uo_out[1].n0 uo_out[1].t3 211.01
R1348 uo_out[1].n1 uo_out[1].n0 152
R1349 uo_out[1].n5 uo_out[1] 12.6752
R1350 uo_out[1].n4 uo_out[1].n1 11.6411
R1351 uo_out[1].n4 uo_out[1].n3 9.3005
R1352 uo_out[1].n3 uo_out[1] 7.17626
R1353 uo_out[1].n3 uo_out[1].n2 4.84898
R1354 uo_out[1].n5 uo_out[1].n4 4.5029
R1355 uo_out[1].n1 uo_out[1] 1.37896
R1356 uo_out[1] uo_out[1].n5 0.0730806
R1357 uo_out[0].n4 uo_out[0].t0 983.422
R1358 uo_out[0] uo_out[0].t1 455.764
R1359 uo_out[0].n0 uo_out[0].t2 294.557
R1360 uo_out[0].n0 uo_out[0].t3 211.01
R1361 uo_out[0].n1 uo_out[0].n0 152
R1362 uo_out[0].n4 uo_out[0].n3 19.6603
R1363 uo_out[0].n2 uo_out[0].n1 17.6405
R1364 uo_out[0] uo_out[0].n4 10.2862
R1365 uo_out[0].n3 uo_out[0].n2 6.83545
R1366 uo_out[0].n1 uo_out[0] 2.01193
R1367 uo_out[0].n3 uo_out[0] 1.31337
R1368 uo_out[0].n2 uo_out[0] 0.0793043
R1369 uo_out[3].n0 uo_out[3].t0 313.104
R1370 uo_out[3].t1 uo_out[3].n0 265.769
R1371 uo_out[3] uo_out[3].t1 262.318
R1372 uo_out[3].n2 uo_out[3] 19.5328
R1373 uo_out[3].n2 uo_out[3].n1 13.8005
R1374 uo_out[3].n1 uo_out[3].n0 7.17626
R1375 uo_out[3].n1 uo_out[3] 4.84898
R1376 uo_out[3] uo_out[3].n2 0.0529194
C0 m2_6582_13386# m1_6582_13386# 2.03601f
C1 m3_12074_25760# m2_12074_25760# 98.466896f
C2 m1_25292_15258# m2_25292_15258# 2.03601f
C3 m1_19762_10378# m2_19762_10378# 2.03601f
C4 m1_13228_33714# m2_13228_33714# 2.03601f
C5 m2_7102_32098# m1_7102_32098# 2.03601f
C6 m2_4034_22148# m1_4034_22148# 2.03601f
C7 m2_3514_25724# m1_3514_25724# 2.03601f
C8 m1_6582_15306# m2_6582_15306# 2.03601f
C9 m2_4568_16810# m1_4568_16810# 2.03601f
C10 m1_16274_9582# m2_16274_9582# 2.03601f
C11 m2_9378_11156# m1_9378_11156# 2.03601f
C12 m1_13228_35634# m2_13228_35634# 2.03601f
C13 m2_7102_30178# m1_7102_30178# 2.03601f
C14 m1_25292_17178# m2_25292_17178# 2.03601f
C15 m2_3514_23804# m1_3514_23804# 2.03601f
C16 m2_25812_28774# m1_25812_28774# 2.03601f
C17 m2_23378_31396# m1_23378_31396# 2.03601f
C18 m2_16794_33982# m1_16794_33982# 2.03601f
C19 m2_16794_35902# m1_16794_35902# 2.03601f
C20 m2_9378_13076# m1_9378_13076# 2.03601f
C21 m2_19762_12298# m1_19762_12298# 2.03601f
C22 m1_22858_12168# m2_22858_12168# 2.03601f
C23 m2_23378_33316# m1_23378_33316# 2.03601f
C24 m1_10514_15880# m2_10514_15880# 0.104063p
C25 m4_12074_25760# m3_12074_25760# 95.99921f
C26 m1_9900_34328# m2_9900_34328# 2.03601f
C27 m1_12708_9850# m2_12708_9850# 2.03601f
C28 m2_20282_35106# m1_20282_35106# 2.03601f
C29 m1_10716_42050# m2_10716_42050# 2.03601f
C30 m2_26844_18480# m1_26844_18480# 2.03601f
C31 m2_4568_18730# m1_4568_18730# 2.03601f
C32 m2_27898_22016# m1_27898_22016# 2.03601f
C33 m2_26844_27472# m1_26844_27472# 2.03601f
C34 m2_5088_27222# m1_5088_27222# 2.03601f
C35 m2_26844_25552# m1_26844_25552# 2.03601f
C36 m1_22858_14088# m2_22858_14088# 2.03601f
C37 m2_5088_29142# m1_5088_29142# 2.03601f
C38 m2_10514_15880# m3_10514_15880# 67.004105f
C39 VAPWR VDPWR 19.2978f
C40 m2_12456_42110# m1_12456_42110# 2.03601f
C41 m1_25812_30694# m2_25812_30694# 2.03601f
C42 m1_16274_11502# m2_16274_11502# 2.03601f
C43 m1_26844_20400# m2_26844_20400# 2.03601f
C44 m1_4034_20228# m2_4034_20228# 2.03601f
C45 m1_27898_23936# m2_27898_23936# 2.03601f
C46 m2_12708_11770# m1_12708_11770# 2.03601f
C47 m4_10514_15880# m3_10514_15880# 65.3249f
C48 m1_9900_32408# m2_9900_32408# 2.03601f
C49 m2_20282_33186# m1_20282_33186# 2.03601f
C50 uo_out[0] VDPWR 2.35179f
C51 m1_12074_25760# m2_12074_25760# 0.152927p
C52 uo_out[0] VGND 4.703662f
C53 uo_out[3] VGND 2.04563f
C54 VAPWR VGND 0.145745p
C55 VDPWR VGND 54.020542f
C56 m4_10514_15880# VGND 11.069901f $ **FLOATING
C57 m4_12074_25760# VGND 8.74745f $ **FLOATING
C58 m3_10514_15880# VGND 12.5706f $ **FLOATING
C59 m3_12074_25760# VGND 10.2013f $ **FLOATING
C60 m2_10514_15880# VGND 11.5361f $ **FLOATING
C61 m2_12074_25760# VGND 9.56453f $ **FLOATING
C62 m1_10514_15880# VGND 32.9027f $ **FLOATING
C63 m1_12074_25760# VGND 40.2807f $ **FLOATING
C64 ring_0/skullfet_inverter_16.A VGND 4.98713f
C65 ring_0/skullfet_inverter_17.A VGND 5.087f
C66 ring_0/skullfet_inverter_15.A VGND 5.26433f
C67 ring_0/skullfet_inverter_18.A VGND 5.29181f
C68 ring_0/skullfet_inverter_14.A VGND 5.42234f
C69 ring_0/skullfet_inverter_19.A VGND 5.55224f
C70 ring_0/skullfet_inverter_13.A VGND 5.39855f
C71 ring_0/skullfet_inverter_20.A VGND 5.37944f
C72 ring_0/skullfet_inverter_12.A VGND 5.705f
C73 ring_0/skullfet_inverter_20.Y VGND 6.09239f
C74 ring_0/skullfet_inverter_11.A VGND 5.64345f
C75 ring_0/skullfet_inverter_1.A VGND 5.89097f
C76 ring_0/skullfet_inverter_10.A VGND 6.07373f
C77 ring_0/skullfet_inverter_2.A VGND 5.83825f
C78 ring_0/skullfet_inverter_9.A VGND 5.19847f
C79 ring_0/skullfet_inverter_3.A VGND 5.40935f
C80 ring_0/skullfet_inverter_4.A VGND 5.35941f
C81 ring_0/skullfet_inverter_8.A VGND 5.38592f
C82 ring_0/skullfet_inverter_6.A VGND 4.983f
C83 ring_0/skullfet_inverter_5.A VGND 5.14674f
C84 skullfet_level_shifter.A VGND 11.6428f
C85 VDPWR.n3 VGND 7.59376f
C86 VAPWR.n103 VGND 2.52536f
C87 VAPWR.n104 VGND 14.571099f
.ends

