VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_oscillating_bones
  CLASS BLOCK ;
  FOREIGN tt_um_oscillating_bones ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 15.434999 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 124.754196 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.000 5.000 6.500 220.760 ;
    END
  END VAPWR
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3.000 5.000 4.500 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 62.600 219.685 91.040 221.290 ;
      LAYER pwell ;
        RECT 62.795 219.165 65.560 219.395 ;
        RECT 67.100 219.165 68.010 219.385 ;
        RECT 62.795 218.485 71.525 219.165 ;
        RECT 71.545 218.570 71.975 219.355 ;
        RECT 72.005 218.570 72.435 219.355 ;
        RECT 72.455 219.165 75.220 219.395 ;
        RECT 76.760 219.165 77.670 219.385 ;
        RECT 72.455 218.485 81.185 219.165 ;
        RECT 81.205 218.570 81.635 219.355 ;
        RECT 81.665 218.570 82.095 219.355 ;
        RECT 82.115 219.165 84.880 219.395 ;
        RECT 86.420 219.165 87.330 219.385 ;
        RECT 82.115 218.485 90.845 219.165 ;
        RECT 71.215 218.295 71.385 218.485 ;
        RECT 80.875 218.295 81.045 218.485 ;
        RECT 90.535 218.295 90.705 218.485 ;
        RECT 53.210 208.740 58.930 214.520 ;
      LAYER nwell ;
        RECT 61.650 208.740 67.990 214.520 ;
      LAYER pwell ;
        RECT 65.470 175.820 71.250 181.540 ;
        RECT 83.300 177.160 89.080 182.880 ;
        RECT 48.830 169.290 54.610 175.010 ;
      LAYER nwell ;
        RECT 65.470 166.760 71.250 173.100 ;
        RECT 83.300 168.100 89.080 174.440 ;
      LAYER pwell ;
        RECT 100.740 173.180 106.520 178.900 ;
        RECT 34.840 158.140 40.620 163.860 ;
      LAYER nwell ;
        RECT 48.830 160.230 54.610 166.570 ;
        RECT 100.740 164.120 106.520 170.460 ;
      LAYER pwell ;
        RECT 116.220 164.230 122.000 169.950 ;
      LAYER nwell ;
        RECT 34.840 149.080 40.620 155.420 ;
        RECT 116.220 155.170 122.000 161.510 ;
      LAYER pwell ;
        RECT 128.390 151.120 134.170 156.840 ;
        RECT 24.770 143.360 30.550 149.080 ;
      LAYER nwell ;
        RECT 128.390 142.060 134.170 148.400 ;
        RECT 24.770 134.300 30.550 140.640 ;
      LAYER pwell ;
        RECT 133.610 135.010 139.390 140.730 ;
        RECT 16.960 126.270 22.740 131.990 ;
      LAYER nwell ;
        RECT 133.610 125.950 139.390 132.290 ;
        RECT 16.960 117.210 22.740 123.550 ;
      LAYER pwell ;
        RECT 138.820 117.330 144.600 123.050 ;
        RECT 19.500 108.390 25.280 114.110 ;
      LAYER nwell ;
        RECT 138.820 108.270 144.600 114.610 ;
        RECT 19.500 99.330 25.280 105.670 ;
      LAYER pwell ;
        RECT 133.610 99.650 139.390 105.370 ;
        RECT 22.230 91.300 28.010 97.020 ;
      LAYER nwell ;
        RECT 133.610 90.590 139.390 96.930 ;
        RECT 22.230 82.240 28.010 88.580 ;
      LAYER pwell ;
        RECT 125.850 83.540 131.630 89.260 ;
      LAYER nwell ;
        RECT 32.300 73.800 38.080 80.140 ;
        RECT 125.850 74.480 131.630 80.820 ;
      LAYER pwell ;
        RECT 32.300 65.360 38.080 71.080 ;
      LAYER nwell ;
        RECT 46.280 62.650 52.060 68.990 ;
        RECT 113.680 67.710 119.460 74.050 ;
      LAYER pwell ;
        RECT 46.280 54.210 52.060 59.930 ;
      LAYER nwell ;
        RECT 62.930 56.120 68.710 62.460 ;
        RECT 80.760 54.780 86.540 61.120 ;
        RECT 98.200 58.760 103.980 65.100 ;
      LAYER pwell ;
        RECT 113.680 59.270 119.460 64.990 ;
        RECT 62.930 47.680 68.710 53.400 ;
        RECT 80.760 46.340 86.540 52.060 ;
        RECT 98.200 50.320 103.980 56.040 ;
      LAYER li1 ;
        RECT 62.790 221.015 90.850 221.185 ;
        RECT 62.880 219.860 63.215 220.845 ;
        RECT 63.385 219.875 63.600 221.015 ;
        RECT 63.790 220.095 64.120 220.825 ;
        RECT 62.880 219.290 63.115 219.860 ;
        RECT 63.790 219.705 64.060 220.095 ;
        RECT 64.310 219.955 64.640 220.800 ;
        RECT 64.810 220.005 64.980 221.015 ;
        RECT 65.150 220.285 65.490 220.845 ;
        RECT 65.725 220.515 66.040 221.015 ;
        RECT 66.220 220.545 67.105 220.715 ;
        RECT 63.285 219.375 64.060 219.705 ;
        RECT 62.880 218.635 63.135 219.290 ;
        RECT 63.860 218.995 64.060 219.375 ;
        RECT 64.230 219.875 64.640 219.955 ;
        RECT 65.150 219.910 66.050 220.285 ;
        RECT 64.230 219.825 64.465 219.875 ;
        RECT 64.230 219.245 64.420 219.825 ;
        RECT 65.150 219.705 65.340 219.910 ;
        RECT 66.220 219.705 66.390 220.545 ;
        RECT 67.330 220.515 67.580 220.845 ;
        RECT 64.590 219.375 65.340 219.705 ;
        RECT 65.510 219.375 66.390 219.705 ;
        RECT 64.230 219.205 64.475 219.245 ;
        RECT 65.140 219.205 65.340 219.375 ;
        RECT 64.230 219.120 64.630 219.205 ;
        RECT 63.305 218.465 63.625 218.925 ;
        RECT 63.860 218.725 64.110 218.995 ;
        RECT 64.300 218.685 64.630 219.120 ;
        RECT 64.800 218.465 64.970 219.075 ;
        RECT 65.140 218.680 65.470 219.205 ;
        RECT 65.735 218.465 65.945 218.995 ;
        RECT 66.220 218.915 66.390 219.375 ;
        RECT 66.560 219.415 66.880 220.375 ;
        RECT 67.050 219.625 67.240 220.345 ;
        RECT 67.410 219.445 67.580 220.515 ;
        RECT 67.750 220.215 67.920 221.015 ;
        RECT 68.090 220.570 69.195 220.740 ;
        RECT 68.090 219.955 68.260 220.570 ;
        RECT 69.405 220.420 69.655 220.845 ;
        RECT 69.825 220.555 70.090 221.015 ;
        RECT 68.430 220.035 68.960 220.400 ;
        RECT 69.405 220.290 69.710 220.420 ;
        RECT 67.750 219.865 68.260 219.955 ;
        RECT 67.750 219.695 68.620 219.865 ;
        RECT 67.750 219.625 67.920 219.695 ;
        RECT 68.040 219.445 68.240 219.475 ;
        RECT 66.560 219.085 67.025 219.415 ;
        RECT 67.410 219.145 68.240 219.445 ;
        RECT 67.410 218.915 67.580 219.145 ;
        RECT 66.220 218.745 67.005 218.915 ;
        RECT 67.175 218.745 67.580 218.915 ;
        RECT 67.760 218.465 68.130 218.965 ;
        RECT 68.450 218.915 68.620 219.695 ;
        RECT 68.790 219.335 68.960 220.035 ;
        RECT 69.130 219.505 69.370 220.100 ;
        RECT 68.790 219.115 69.315 219.335 ;
        RECT 69.540 219.185 69.710 220.290 ;
        RECT 69.485 219.055 69.710 219.185 ;
        RECT 69.880 219.095 70.160 220.045 ;
        RECT 69.485 218.915 69.655 219.055 ;
        RECT 68.450 218.745 69.125 218.915 ;
        RECT 69.320 218.745 69.655 218.915 ;
        RECT 69.825 218.465 70.075 218.925 ;
        RECT 70.330 218.725 70.515 220.845 ;
        RECT 70.685 220.515 71.015 221.015 ;
        RECT 71.185 220.345 71.355 220.845 ;
        RECT 70.690 220.175 71.355 220.345 ;
        RECT 70.690 219.185 70.920 220.175 ;
        RECT 71.090 219.355 71.440 220.005 ;
        RECT 71.615 219.850 71.905 221.015 ;
        RECT 72.075 219.850 72.365 221.015 ;
        RECT 72.540 219.860 72.875 220.845 ;
        RECT 73.045 219.875 73.260 221.015 ;
        RECT 73.450 220.095 73.780 220.825 ;
        RECT 72.540 219.290 72.775 219.860 ;
        RECT 73.450 219.705 73.720 220.095 ;
        RECT 73.970 219.955 74.300 220.800 ;
        RECT 74.470 220.005 74.640 221.015 ;
        RECT 74.810 220.285 75.150 220.845 ;
        RECT 75.385 220.515 75.700 221.015 ;
        RECT 75.880 220.545 76.765 220.715 ;
        RECT 72.945 219.375 73.720 219.705 ;
        RECT 70.690 219.015 71.355 219.185 ;
        RECT 70.685 218.465 71.015 218.845 ;
        RECT 71.185 218.725 71.355 219.015 ;
        RECT 71.615 218.465 71.905 219.190 ;
        RECT 72.075 218.465 72.365 219.190 ;
        RECT 72.540 218.635 72.795 219.290 ;
        RECT 73.520 218.995 73.720 219.375 ;
        RECT 73.890 219.875 74.300 219.955 ;
        RECT 74.810 219.910 75.710 220.285 ;
        RECT 73.890 219.825 74.125 219.875 ;
        RECT 73.890 219.245 74.080 219.825 ;
        RECT 74.810 219.705 75.000 219.910 ;
        RECT 75.880 219.705 76.050 220.545 ;
        RECT 76.990 220.515 77.240 220.845 ;
        RECT 74.250 219.375 75.000 219.705 ;
        RECT 75.170 219.375 76.050 219.705 ;
        RECT 73.890 219.205 74.135 219.245 ;
        RECT 74.800 219.205 75.000 219.375 ;
        RECT 73.890 219.120 74.290 219.205 ;
        RECT 72.965 218.465 73.285 218.925 ;
        RECT 73.520 218.725 73.770 218.995 ;
        RECT 73.960 218.685 74.290 219.120 ;
        RECT 74.460 218.465 74.630 219.075 ;
        RECT 74.800 218.680 75.130 219.205 ;
        RECT 75.395 218.465 75.605 218.995 ;
        RECT 75.880 218.915 76.050 219.375 ;
        RECT 76.220 219.415 76.540 220.375 ;
        RECT 76.710 219.625 76.900 220.345 ;
        RECT 77.070 219.445 77.240 220.515 ;
        RECT 77.410 220.215 77.580 221.015 ;
        RECT 77.750 220.570 78.855 220.740 ;
        RECT 77.750 219.955 77.920 220.570 ;
        RECT 79.065 220.420 79.315 220.845 ;
        RECT 79.485 220.555 79.750 221.015 ;
        RECT 78.090 220.035 78.620 220.400 ;
        RECT 79.065 220.290 79.370 220.420 ;
        RECT 77.410 219.865 77.920 219.955 ;
        RECT 77.410 219.695 78.280 219.865 ;
        RECT 77.410 219.625 77.580 219.695 ;
        RECT 77.700 219.445 77.900 219.475 ;
        RECT 76.220 219.085 76.685 219.415 ;
        RECT 77.070 219.145 77.900 219.445 ;
        RECT 77.070 218.915 77.240 219.145 ;
        RECT 75.880 218.745 76.665 218.915 ;
        RECT 76.835 218.745 77.240 218.915 ;
        RECT 77.420 218.465 77.790 218.965 ;
        RECT 78.110 218.915 78.280 219.695 ;
        RECT 78.450 219.335 78.620 220.035 ;
        RECT 78.790 219.505 79.030 220.100 ;
        RECT 78.450 219.115 78.975 219.335 ;
        RECT 79.200 219.185 79.370 220.290 ;
        RECT 79.145 219.055 79.370 219.185 ;
        RECT 79.540 219.095 79.820 220.045 ;
        RECT 79.145 218.915 79.315 219.055 ;
        RECT 78.110 218.745 78.785 218.915 ;
        RECT 78.980 218.745 79.315 218.915 ;
        RECT 79.485 218.465 79.735 218.925 ;
        RECT 79.990 218.725 80.175 220.845 ;
        RECT 80.345 220.515 80.675 221.015 ;
        RECT 80.845 220.345 81.015 220.845 ;
        RECT 80.350 220.175 81.015 220.345 ;
        RECT 80.350 219.185 80.580 220.175 ;
        RECT 80.750 219.355 81.100 220.005 ;
        RECT 81.275 219.850 81.565 221.015 ;
        RECT 81.735 219.850 82.025 221.015 ;
        RECT 82.200 219.860 82.535 220.845 ;
        RECT 82.705 219.875 82.920 221.015 ;
        RECT 83.110 220.095 83.440 220.825 ;
        RECT 82.200 219.290 82.435 219.860 ;
        RECT 83.110 219.705 83.380 220.095 ;
        RECT 83.630 219.955 83.960 220.800 ;
        RECT 84.130 220.005 84.300 221.015 ;
        RECT 84.470 220.285 84.810 220.845 ;
        RECT 85.045 220.515 85.360 221.015 ;
        RECT 85.540 220.545 86.425 220.715 ;
        RECT 82.605 219.375 83.380 219.705 ;
        RECT 80.350 219.015 81.015 219.185 ;
        RECT 80.345 218.465 80.675 218.845 ;
        RECT 80.845 218.725 81.015 219.015 ;
        RECT 81.275 218.465 81.565 219.190 ;
        RECT 81.735 218.465 82.025 219.190 ;
        RECT 82.200 218.635 82.455 219.290 ;
        RECT 83.180 218.995 83.380 219.375 ;
        RECT 83.550 219.875 83.960 219.955 ;
        RECT 84.470 219.910 85.370 220.285 ;
        RECT 83.550 219.825 83.785 219.875 ;
        RECT 83.550 219.245 83.740 219.825 ;
        RECT 84.470 219.705 84.660 219.910 ;
        RECT 85.540 219.705 85.710 220.545 ;
        RECT 86.650 220.515 86.900 220.845 ;
        RECT 83.910 219.375 84.660 219.705 ;
        RECT 84.830 219.375 85.710 219.705 ;
        RECT 83.550 219.205 83.795 219.245 ;
        RECT 84.460 219.205 84.660 219.375 ;
        RECT 83.550 219.120 83.950 219.205 ;
        RECT 82.625 218.465 82.945 218.925 ;
        RECT 83.180 218.725 83.430 218.995 ;
        RECT 83.620 218.685 83.950 219.120 ;
        RECT 84.120 218.465 84.290 219.075 ;
        RECT 84.460 218.680 84.790 219.205 ;
        RECT 85.055 218.465 85.265 218.995 ;
        RECT 85.540 218.915 85.710 219.375 ;
        RECT 85.880 219.415 86.200 220.375 ;
        RECT 86.370 219.625 86.560 220.345 ;
        RECT 86.730 219.445 86.900 220.515 ;
        RECT 87.070 220.215 87.240 221.015 ;
        RECT 87.410 220.570 88.515 220.740 ;
        RECT 87.410 219.955 87.580 220.570 ;
        RECT 88.725 220.420 88.975 220.845 ;
        RECT 89.145 220.555 89.410 221.015 ;
        RECT 87.750 220.035 88.280 220.400 ;
        RECT 88.725 220.290 89.030 220.420 ;
        RECT 87.070 219.865 87.580 219.955 ;
        RECT 87.070 219.695 87.940 219.865 ;
        RECT 87.070 219.625 87.240 219.695 ;
        RECT 87.360 219.445 87.560 219.475 ;
        RECT 85.880 219.085 86.345 219.415 ;
        RECT 86.730 219.145 87.560 219.445 ;
        RECT 86.730 218.915 86.900 219.145 ;
        RECT 85.540 218.745 86.325 218.915 ;
        RECT 86.495 218.745 86.900 218.915 ;
        RECT 87.080 218.465 87.450 218.965 ;
        RECT 87.770 218.915 87.940 219.695 ;
        RECT 88.110 219.335 88.280 220.035 ;
        RECT 88.450 219.505 88.690 220.100 ;
        RECT 88.110 219.115 88.635 219.335 ;
        RECT 88.860 219.185 89.030 220.290 ;
        RECT 88.805 219.055 89.030 219.185 ;
        RECT 89.200 219.095 89.480 220.045 ;
        RECT 88.805 218.915 88.975 219.055 ;
        RECT 87.770 218.745 88.445 218.915 ;
        RECT 88.640 218.745 88.975 218.915 ;
        RECT 89.145 218.465 89.395 218.925 ;
        RECT 89.650 218.725 89.835 220.845 ;
        RECT 90.005 220.515 90.335 221.015 ;
        RECT 90.505 220.345 90.675 220.845 ;
        RECT 90.010 220.175 90.675 220.345 ;
        RECT 90.010 219.185 90.240 220.175 ;
        RECT 90.410 219.355 90.760 220.005 ;
        RECT 90.010 219.015 90.675 219.185 ;
        RECT 90.005 218.465 90.335 218.845 ;
        RECT 90.505 218.725 90.675 219.015 ;
        RECT 62.790 218.295 90.850 218.465 ;
        RECT 55.710 214.570 65.270 215.130 ;
        RECT 54.150 214.240 54.710 214.460 ;
        RECT 53.320 213.350 54.710 214.240 ;
        RECT 55.710 213.460 56.270 214.570 ;
        RECT 64.710 213.350 65.270 214.570 ;
        RECT 66.820 214.130 67.600 214.180 ;
        RECT 66.270 213.400 67.600 214.130 ;
        RECT 54.150 213.130 54.710 213.350 ;
        RECT 66.270 213.130 66.820 213.400 ;
        RECT 57.600 207.900 63.600 208.460 ;
        RECT 83.580 181.940 84.470 182.770 ;
        RECT 65.750 180.600 66.640 181.430 ;
        RECT 83.360 181.380 84.690 181.940 ;
        RECT 65.530 180.040 66.860 180.600 ;
        RECT 82.690 179.820 84.360 180.380 ;
        RECT 64.860 178.480 66.530 179.040 ;
        RECT 49.110 174.070 50.000 174.900 ;
        RECT 48.890 173.510 50.220 174.070 ;
        RECT 48.220 171.950 49.890 172.510 ;
        RECT 35.120 162.920 36.010 163.750 ;
        RECT 48.220 163.510 48.780 171.950 ;
        RECT 54.890 164.620 55.450 170.620 ;
        RECT 64.860 170.040 65.420 178.480 ;
        RECT 71.530 171.150 72.090 177.150 ;
        RECT 82.690 171.380 83.250 179.820 ;
        RECT 89.360 172.490 89.920 178.490 ;
        RECT 101.020 177.960 101.910 178.790 ;
        RECT 100.800 177.400 102.130 177.960 ;
        RECT 100.130 175.840 101.800 176.400 ;
        RECT 82.690 170.820 84.470 171.380 ;
        RECT 64.860 169.480 66.640 170.040 ;
        RECT 83.690 169.270 84.690 169.820 ;
        RECT 83.640 168.490 84.420 169.270 ;
        RECT 65.860 167.930 66.860 168.480 ;
        RECT 65.810 167.150 66.590 167.930 ;
        RECT 100.130 167.400 100.690 175.840 ;
        RECT 106.800 168.510 107.360 174.510 ;
        RECT 116.500 169.010 117.390 169.840 ;
        RECT 116.280 168.450 117.610 169.010 ;
        RECT 100.130 166.840 101.910 167.400 ;
        RECT 115.610 166.890 117.280 167.450 ;
        RECT 101.130 165.290 102.130 165.840 ;
        RECT 101.080 164.510 101.860 165.290 ;
        RECT 48.220 162.950 50.000 163.510 ;
        RECT 34.900 162.360 36.230 162.920 ;
        RECT 49.220 161.400 50.220 161.950 ;
        RECT 34.230 160.800 35.900 161.360 ;
        RECT 34.230 152.360 34.790 160.800 ;
        RECT 49.170 160.620 49.950 161.400 ;
        RECT 40.900 153.470 41.460 159.470 ;
        RECT 115.610 158.450 116.170 166.890 ;
        RECT 122.280 159.560 122.840 165.560 ;
        RECT 115.610 157.890 117.390 158.450 ;
        RECT 116.610 156.340 117.610 156.890 ;
        RECT 116.560 155.560 117.340 156.340 ;
        RECT 128.670 155.900 129.560 156.730 ;
        RECT 128.450 155.340 129.780 155.900 ;
        RECT 127.780 153.780 129.450 154.340 ;
        RECT 34.230 151.800 36.010 152.360 ;
        RECT 35.230 150.250 36.230 150.800 ;
        RECT 35.180 149.470 35.960 150.250 ;
        RECT 25.050 148.140 25.940 148.970 ;
        RECT 24.830 147.580 26.160 148.140 ;
        RECT 24.160 146.020 25.830 146.580 ;
        RECT 24.160 137.580 24.720 146.020 ;
        RECT 127.780 145.340 128.340 153.780 ;
        RECT 134.450 146.450 135.010 152.450 ;
        RECT 127.780 144.780 129.560 145.340 ;
        RECT 30.830 138.690 31.390 144.690 ;
        RECT 128.780 143.230 129.780 143.780 ;
        RECT 128.730 142.450 129.510 143.230 ;
        RECT 138.220 139.790 139.110 140.620 ;
        RECT 138.000 139.230 139.330 139.790 ;
        RECT 138.330 137.670 140.000 138.230 ;
        RECT 24.160 137.020 25.940 137.580 ;
        RECT 25.160 135.470 26.160 136.020 ;
        RECT 25.110 134.690 25.890 135.470 ;
        RECT 21.570 131.050 22.460 131.880 ;
        RECT 21.350 130.490 22.680 131.050 ;
        RECT 132.770 130.340 133.330 136.340 ;
        RECT 21.680 128.930 23.350 129.490 ;
        RECT 139.440 129.230 140.000 137.670 ;
        RECT 16.120 121.600 16.680 127.600 ;
        RECT 22.790 120.490 23.350 128.930 ;
        RECT 138.220 128.670 140.000 129.230 ;
        RECT 138.000 127.120 139.000 127.670 ;
        RECT 138.270 126.340 139.050 127.120 ;
        RECT 139.100 122.110 139.990 122.940 ;
        RECT 138.880 121.550 140.210 122.110 ;
        RECT 21.570 119.930 23.350 120.490 ;
        RECT 138.210 119.990 139.880 120.550 ;
        RECT 21.350 118.380 22.350 118.930 ;
        RECT 21.620 117.600 22.400 118.380 ;
        RECT 19.780 113.170 20.670 114.000 ;
        RECT 19.560 112.610 20.890 113.170 ;
        RECT 18.890 111.050 20.560 111.610 ;
        RECT 138.210 111.550 138.770 119.990 ;
        RECT 144.880 112.660 145.440 118.660 ;
        RECT 18.890 102.610 19.450 111.050 ;
        RECT 138.210 110.990 139.990 111.550 ;
        RECT 25.560 103.720 26.120 109.720 ;
        RECT 139.210 109.440 140.210 109.990 ;
        RECT 139.160 108.660 139.940 109.440 ;
        RECT 138.220 104.430 139.110 105.260 ;
        RECT 138.000 103.870 139.330 104.430 ;
        RECT 18.890 102.050 20.670 102.610 ;
        RECT 138.330 102.310 140.000 102.870 ;
        RECT 19.890 100.500 20.890 101.050 ;
        RECT 19.840 99.720 20.620 100.500 ;
        RECT 26.840 96.080 27.730 96.910 ;
        RECT 26.620 95.520 27.950 96.080 ;
        RECT 132.770 94.980 133.330 100.980 ;
        RECT 26.950 93.960 28.620 94.520 ;
        RECT 21.390 86.630 21.950 92.630 ;
        RECT 28.060 85.520 28.620 93.960 ;
        RECT 139.440 93.870 140.000 102.310 ;
        RECT 138.220 93.310 140.000 93.870 ;
        RECT 138.000 91.760 139.000 92.310 ;
        RECT 138.270 90.980 139.050 91.760 ;
        RECT 130.460 88.320 131.350 89.150 ;
        RECT 130.240 87.760 131.570 88.320 ;
        RECT 130.570 86.200 132.240 86.760 ;
        RECT 26.840 84.960 28.620 85.520 ;
        RECT 26.620 83.410 27.620 83.960 ;
        RECT 26.890 82.630 27.670 83.410 ;
        RECT 36.960 78.970 37.740 79.750 ;
        RECT 36.690 78.420 37.690 78.970 ;
        RECT 125.010 78.870 125.570 84.870 ;
        RECT 131.680 77.760 132.240 86.200 ;
        RECT 36.910 76.860 38.690 77.420 ;
        RECT 130.460 77.200 132.240 77.760 ;
        RECT 31.460 69.750 32.020 75.750 ;
        RECT 38.130 68.420 38.690 76.860 ;
        RECT 130.240 75.650 131.240 76.200 ;
        RECT 130.510 74.870 131.290 75.650 ;
        RECT 118.340 72.880 119.120 73.660 ;
        RECT 118.070 72.330 119.070 72.880 ;
        RECT 118.290 70.770 120.070 71.330 ;
        RECT 37.020 67.860 38.690 68.420 ;
        RECT 50.940 67.820 51.720 68.600 ;
        RECT 50.670 67.270 51.670 67.820 ;
        RECT 36.690 66.300 38.020 66.860 ;
        RECT 36.910 65.470 37.800 66.300 ;
        RECT 50.890 65.710 52.670 66.270 ;
        RECT 45.440 58.600 46.000 64.600 ;
        RECT 52.110 57.270 52.670 65.710 ;
        RECT 102.860 63.930 103.640 64.710 ;
        RECT 102.590 63.380 103.590 63.930 ;
        RECT 112.840 63.660 113.400 69.660 ;
        RECT 67.590 61.290 68.370 62.070 ;
        RECT 102.810 61.820 104.590 62.380 ;
        RECT 119.510 62.330 120.070 70.770 ;
        RECT 67.320 60.740 68.320 61.290 ;
        RECT 85.420 59.950 86.200 60.730 ;
        RECT 67.540 59.180 69.320 59.740 ;
        RECT 85.150 59.400 86.150 59.950 ;
        RECT 51.000 56.710 52.670 57.270 ;
        RECT 50.670 55.150 52.000 55.710 ;
        RECT 50.890 54.320 51.780 55.150 ;
        RECT 62.090 52.070 62.650 58.070 ;
        RECT 68.760 50.740 69.320 59.180 ;
        RECT 85.370 57.840 87.150 58.400 ;
        RECT 67.650 50.180 69.320 50.740 ;
        RECT 79.920 50.730 80.480 56.730 ;
        RECT 86.590 49.400 87.150 57.840 ;
        RECT 97.360 54.710 97.920 60.710 ;
        RECT 104.030 53.380 104.590 61.820 ;
        RECT 118.400 61.770 120.070 62.330 ;
        RECT 118.070 60.210 119.400 60.770 ;
        RECT 118.290 59.380 119.180 60.210 ;
        RECT 102.920 52.820 104.590 53.380 ;
        RECT 102.590 51.260 103.920 51.820 ;
        RECT 102.810 50.430 103.700 51.260 ;
        RECT 67.320 48.620 68.650 49.180 ;
        RECT 85.480 48.840 87.150 49.400 ;
        RECT 67.540 47.790 68.430 48.620 ;
        RECT 85.150 47.280 86.480 47.840 ;
        RECT 85.370 46.450 86.260 47.280 ;
      LAYER met1 ;
        RECT 90.535 221.340 92.300 221.345 ;
        RECT 62.790 220.865 92.300 221.340 ;
        RECT 62.790 220.860 90.850 220.865 ;
        RECT 67.000 220.320 67.290 220.365 ;
        RECT 68.570 220.320 68.860 220.365 ;
        RECT 70.670 220.320 70.960 220.365 ;
        RECT 67.000 220.180 70.960 220.320 ;
        RECT 67.000 220.135 67.290 220.180 ;
        RECT 68.570 220.135 68.860 220.180 ;
        RECT 70.670 220.135 70.960 220.180 ;
        RECT 76.660 220.320 76.950 220.365 ;
        RECT 78.230 220.320 78.520 220.365 ;
        RECT 80.330 220.320 80.620 220.365 ;
        RECT 76.660 220.180 80.620 220.320 ;
        RECT 76.660 220.135 76.950 220.180 ;
        RECT 78.230 220.135 78.520 220.180 ;
        RECT 80.330 220.135 80.620 220.180 ;
        RECT 86.320 220.320 86.610 220.365 ;
        RECT 87.890 220.320 88.180 220.365 ;
        RECT 89.990 220.320 90.280 220.365 ;
        RECT 86.320 220.180 90.280 220.320 ;
        RECT 86.320 220.135 86.610 220.180 ;
        RECT 87.890 220.135 88.180 220.180 ;
        RECT 89.990 220.135 90.280 220.180 ;
        RECT 62.880 219.870 63.170 220.100 ;
        RECT 66.565 219.980 66.855 220.025 ;
        RECT 69.085 219.980 69.375 220.025 ;
        RECT 70.275 219.980 70.565 220.025 ;
        RECT 62.990 219.640 63.130 219.870 ;
        RECT 66.565 219.840 70.565 219.980 ;
        RECT 72.535 219.870 72.825 220.100 ;
        RECT 76.225 219.980 76.515 220.025 ;
        RECT 78.745 219.980 79.035 220.025 ;
        RECT 79.935 219.980 80.225 220.025 ;
        RECT 66.565 219.795 66.855 219.840 ;
        RECT 69.085 219.795 69.375 219.840 ;
        RECT 70.275 219.795 70.565 219.840 ;
        RECT 69.850 219.640 70.140 219.680 ;
        RECT 62.990 219.500 70.140 219.640 ;
        RECT 69.850 219.450 70.140 219.500 ;
        RECT 71.140 219.425 71.430 219.655 ;
        RECT 72.645 219.640 72.785 219.870 ;
        RECT 76.225 219.840 80.225 219.980 ;
        RECT 82.200 219.870 82.490 220.100 ;
        RECT 85.885 219.980 86.175 220.025 ;
        RECT 88.405 219.980 88.695 220.025 ;
        RECT 89.595 219.980 89.885 220.025 ;
        RECT 76.225 219.795 76.515 219.840 ;
        RECT 78.745 219.795 79.035 219.840 ;
        RECT 79.935 219.795 80.225 219.840 ;
        RECT 79.505 219.640 79.795 219.680 ;
        RECT 72.645 219.500 79.795 219.640 ;
        RECT 79.505 219.450 79.795 219.500 ;
        RECT 80.800 219.425 81.090 219.655 ;
        RECT 82.310 219.640 82.450 219.870 ;
        RECT 85.885 219.840 89.885 219.980 ;
        RECT 90.440 219.840 90.720 219.900 ;
        RECT 85.885 219.795 86.175 219.840 ;
        RECT 88.405 219.795 88.695 219.840 ;
        RECT 89.595 219.795 89.885 219.840 ;
        RECT 89.170 219.640 89.460 219.680 ;
        RECT 82.310 219.500 89.460 219.640 ;
        RECT 89.170 219.450 89.460 219.500 ;
        RECT 90.380 219.455 90.740 219.840 ;
        RECT 64.260 218.770 64.690 219.090 ;
        RECT 71.200 219.075 71.370 219.425 ;
        RECT 73.975 219.075 74.265 219.105 ;
        RECT 71.200 219.020 74.265 219.075 ;
        RECT 80.860 219.075 81.030 219.425 ;
        RECT 90.440 219.395 90.720 219.455 ;
        RECT 83.580 219.075 83.990 219.120 ;
        RECT 71.200 218.905 74.350 219.020 ;
        RECT 80.860 218.905 83.990 219.075 ;
        RECT 73.940 218.760 74.350 218.905 ;
        RECT 83.580 218.860 83.990 218.905 ;
        RECT 61.430 218.140 90.850 218.620 ;
        RECT 67.160 216.130 67.820 216.690 ;
        RECT 60.050 215.630 60.700 215.725 ;
        RECT 52.150 214.685 52.750 215.185 ;
        RECT 54.040 214.680 54.650 215.130 ;
        RECT 54.150 214.020 54.650 214.680 ;
        RECT 58.680 214.450 59.280 214.750 ;
        RECT 59.880 214.570 60.880 215.630 ;
        RECT 61.380 214.450 62.280 214.750 ;
        RECT 66.380 214.570 66.990 215.130 ;
        RECT 54.780 213.550 56.580 213.850 ;
        RECT 58.380 213.550 59.580 214.450 ;
        RECT 61.080 214.150 62.580 214.450 ;
        RECT 61.080 213.850 62.280 214.150 ;
        RECT 61.080 213.550 61.980 213.850 ;
        RECT 64.380 213.550 66.180 213.850 ;
        RECT 66.380 213.740 66.820 214.570 ;
        RECT 54.180 213.250 57.480 213.550 ;
        RECT 58.680 213.250 59.880 213.550 ;
        RECT 54.180 212.950 56.280 213.250 ;
        RECT 56.880 212.950 57.480 213.250 ;
        RECT 59.280 212.950 59.880 213.250 ;
        RECT 61.080 212.950 61.680 213.550 ;
        RECT 63.480 213.250 66.780 213.550 ;
        RECT 63.480 212.950 64.080 213.250 ;
        RECT 64.680 212.950 66.780 213.250 ;
        RECT 53.880 212.650 55.980 212.950 ;
        RECT 53.580 212.050 55.980 212.650 ;
        RECT 57.180 212.650 57.780 212.950 ;
        RECT 59.280 212.650 60.180 212.950 ;
        RECT 57.180 212.350 58.680 212.650 ;
        RECT 59.580 212.350 60.180 212.650 ;
        RECT 60.780 212.350 61.380 212.950 ;
        RECT 63.180 212.650 63.780 212.950 ;
        RECT 62.280 212.350 63.780 212.650 ;
        RECT 64.980 212.650 67.080 212.950 ;
        RECT 56.880 212.050 58.380 212.350 ;
        RECT 53.580 211.750 57.480 212.050 ;
        RECT 57.780 211.750 58.680 212.050 ;
        RECT 59.880 211.750 61.080 212.350 ;
        RECT 62.580 212.050 64.080 212.350 ;
        RECT 64.980 212.050 67.380 212.650 ;
        RECT 62.280 211.750 63.180 212.050 ;
        RECT 63.480 211.750 67.380 212.050 ;
        RECT 53.580 211.450 57.180 211.750 ;
        RECT 57.780 211.450 58.380 211.750 ;
        RECT 60.180 211.450 60.780 211.750 ;
        RECT 62.580 211.450 63.180 211.750 ;
        RECT 63.780 211.450 67.380 211.750 ;
        RECT 53.580 211.150 57.480 211.450 ;
        RECT 57.780 211.150 58.680 211.450 ;
        RECT 53.580 210.250 55.980 211.150 ;
        RECT 56.880 210.850 58.380 211.150 ;
        RECT 59.880 210.850 61.080 211.450 ;
        RECT 62.280 211.150 63.180 211.450 ;
        RECT 63.480 211.150 67.380 211.450 ;
        RECT 62.580 210.850 64.080 211.150 ;
        RECT 57.180 210.550 58.680 210.850 ;
        RECT 59.580 210.550 60.180 210.850 ;
        RECT 57.180 210.250 57.780 210.550 ;
        RECT 54.180 209.950 56.280 210.250 ;
        RECT 56.880 209.950 57.780 210.250 ;
        RECT 59.280 210.250 60.180 210.550 ;
        RECT 60.780 210.250 61.380 210.850 ;
        RECT 62.280 210.550 63.780 210.850 ;
        RECT 63.180 210.250 63.780 210.550 ;
        RECT 64.980 210.250 67.380 211.150 ;
        RECT 59.280 209.950 59.880 210.250 ;
        RECT 54.180 209.650 57.180 209.950 ;
        RECT 58.680 209.650 59.880 209.950 ;
        RECT 61.080 209.650 61.680 210.250 ;
        RECT 63.180 209.950 64.080 210.250 ;
        RECT 64.680 209.950 66.780 210.250 ;
        RECT 63.780 209.650 66.780 209.950 ;
        RECT 54.780 209.350 56.580 209.650 ;
        RECT 58.380 208.750 59.580 209.650 ;
        RECT 61.080 209.350 61.980 209.650 ;
        RECT 64.380 209.350 66.180 209.650 ;
        RECT 61.080 209.050 62.280 209.350 ;
        RECT 61.080 208.750 62.580 209.050 ;
        RECT 58.680 208.450 59.280 208.750 ;
        RECT 59.880 207.350 60.880 208.460 ;
        RECT 61.080 208.450 62.280 208.750 ;
        RECT 50.700 174.340 53.100 174.640 ;
        RECT 48.220 174.070 48.670 174.180 ;
        RECT 48.220 173.570 49.330 174.070 ;
        RECT 50.400 174.040 53.100 174.340 ;
        RECT 60.120 174.610 60.620 207.350 ;
        RECT 85.170 182.210 87.570 182.510 ;
        RECT 82.690 181.940 83.140 182.050 ;
        RECT 82.690 181.440 83.800 181.940 ;
        RECT 84.870 181.910 87.570 182.210 ;
        RECT 84.270 181.310 88.170 181.910 ;
        RECT 67.340 180.870 69.740 181.170 ;
        RECT 64.860 180.600 65.310 180.710 ;
        RECT 64.860 180.100 65.970 180.600 ;
        RECT 67.040 180.570 69.740 180.870 ;
        RECT 66.440 179.970 70.340 180.570 ;
        RECT 83.970 180.110 88.470 181.310 ;
        RECT 66.140 178.770 70.640 179.970 ;
        RECT 83.970 179.810 84.870 180.110 ;
        RECT 83.970 179.510 84.570 179.810 ;
        RECT 66.140 178.470 67.040 178.770 ;
        RECT 66.140 178.170 66.740 178.470 ;
        RECT 66.440 177.870 66.740 178.170 ;
        RECT 67.940 177.870 68.840 178.770 ;
        RECT 69.740 178.470 70.640 178.770 ;
        RECT 84.270 179.210 84.570 179.510 ;
        RECT 85.770 179.210 86.670 180.110 ;
        RECT 87.570 179.810 88.470 180.110 ;
        RECT 87.870 179.510 88.470 179.810 ;
        RECT 87.870 179.210 88.170 179.510 ;
        RECT 84.270 178.910 84.870 179.210 ;
        RECT 85.470 178.910 86.970 179.210 ;
        RECT 87.570 178.910 88.170 179.210 ;
        RECT 84.270 178.610 86.070 178.910 ;
        RECT 86.370 178.610 87.870 178.910 ;
        RECT 70.040 178.170 70.640 178.470 ;
        RECT 84.870 178.310 85.770 178.610 ;
        RECT 86.670 178.310 87.870 178.610 ;
        RECT 70.040 177.870 70.340 178.170 ;
        RECT 66.440 177.570 67.040 177.870 ;
        RECT 67.640 177.570 69.140 177.870 ;
        RECT 69.740 177.570 70.340 177.870 ;
        RECT 85.170 177.710 87.270 178.310 ;
        RECT 102.610 178.230 105.010 178.530 ;
        RECT 100.130 177.960 100.580 178.070 ;
        RECT 66.440 177.270 68.240 177.570 ;
        RECT 68.540 177.270 70.040 177.570 ;
        RECT 83.370 177.410 84.270 177.710 ;
        RECT 85.170 177.410 85.470 177.710 ;
        RECT 85.770 177.410 86.070 177.710 ;
        RECT 86.370 177.410 86.670 177.710 ;
        RECT 86.970 177.410 87.270 177.710 ;
        RECT 88.170 177.410 89.070 177.710 ;
        RECT 100.130 177.460 101.240 177.960 ;
        RECT 102.310 177.930 105.010 178.230 ;
        RECT 67.040 176.970 67.940 177.270 ;
        RECT 68.840 176.970 70.040 177.270 ;
        RECT 67.340 176.370 69.440 176.970 ;
        RECT 83.070 176.810 84.570 177.410 ;
        RECT 87.870 176.810 89.370 177.410 ;
        RECT 101.710 177.330 105.610 177.930 ;
        RECT 83.370 176.510 85.170 176.810 ;
        RECT 87.270 176.510 89.070 176.810 ;
        RECT 65.540 176.070 66.440 176.370 ;
        RECT 67.340 176.070 67.640 176.370 ;
        RECT 67.940 176.070 68.240 176.370 ;
        RECT 68.540 176.070 68.840 176.370 ;
        RECT 69.140 176.070 69.440 176.370 ;
        RECT 70.340 176.070 71.240 176.370 ;
        RECT 84.270 176.210 85.470 176.510 ;
        RECT 86.970 176.210 88.170 176.510 ;
        RECT 65.240 175.470 66.740 176.070 ;
        RECT 70.040 175.470 71.540 176.070 ;
        RECT 82.190 175.940 83.250 176.210 ;
        RECT 65.540 175.170 67.340 175.470 ;
        RECT 69.440 175.170 71.240 175.470 ;
        RECT 76.660 175.440 83.250 175.940 ;
        RECT 84.870 175.910 86.070 176.210 ;
        RECT 86.370 175.910 87.570 176.210 ;
        RECT 89.360 175.940 90.470 176.210 ;
        RECT 101.410 176.130 105.910 177.330 ;
        RECT 66.440 174.870 67.640 175.170 ;
        RECT 69.140 174.870 70.340 175.170 ;
        RECT 60.120 174.600 64.210 174.610 ;
        RECT 64.360 174.600 65.420 174.870 ;
        RECT 60.120 174.110 65.420 174.600 ;
        RECT 67.040 174.570 68.240 174.870 ;
        RECT 68.540 174.570 69.740 174.870 ;
        RECT 71.530 174.600 72.640 174.870 ;
        RECT 76.660 174.600 77.160 175.440 ;
        RECT 82.190 175.210 83.250 175.440 ;
        RECT 85.470 175.310 86.970 175.910 ;
        RECT 89.360 175.440 95.090 175.940 ;
        RECT 101.410 175.830 102.310 176.130 ;
        RECT 101.410 175.530 102.010 175.830 ;
        RECT 84.870 175.010 86.070 175.310 ;
        RECT 86.370 175.010 87.570 175.310 ;
        RECT 89.360 175.210 90.470 175.440 ;
        RECT 83.370 174.710 85.470 175.010 ;
        RECT 86.970 174.710 89.370 175.010 ;
        RECT 49.800 173.440 53.700 174.040 ;
        RECT 49.500 172.240 54.000 173.440 ;
        RECT 49.500 171.940 50.400 172.240 ;
        RECT 49.500 171.640 50.100 171.940 ;
        RECT 49.800 171.340 50.100 171.640 ;
        RECT 51.300 171.340 52.200 172.240 ;
        RECT 53.100 171.940 54.000 172.240 ;
        RECT 53.400 171.640 54.000 171.940 ;
        RECT 53.400 171.340 53.700 171.640 ;
        RECT 49.800 171.040 50.400 171.340 ;
        RECT 51.000 171.040 52.500 171.340 ;
        RECT 53.100 171.040 53.700 171.340 ;
        RECT 49.800 170.740 51.600 171.040 ;
        RECT 51.900 170.740 53.400 171.040 ;
        RECT 50.400 170.440 51.300 170.740 ;
        RECT 52.200 170.440 53.400 170.740 ;
        RECT 50.700 169.840 52.800 170.440 ;
        RECT 48.900 169.540 49.800 169.840 ;
        RECT 50.700 169.540 51.000 169.840 ;
        RECT 51.300 169.540 51.600 169.840 ;
        RECT 51.900 169.540 52.200 169.840 ;
        RECT 52.500 169.540 52.800 169.840 ;
        RECT 53.700 169.540 54.600 169.840 ;
        RECT 48.600 168.940 50.100 169.540 ;
        RECT 53.400 168.940 54.900 169.540 ;
        RECT 48.900 168.640 50.700 168.940 ;
        RECT 52.800 168.640 54.600 168.940 ;
        RECT 49.800 168.340 51.000 168.640 ;
        RECT 52.500 168.340 53.700 168.640 ;
        RECT 44.210 168.070 47.580 168.090 ;
        RECT 47.720 168.070 48.780 168.340 ;
        RECT 44.210 167.590 48.780 168.070 ;
        RECT 50.400 168.040 51.600 168.340 ;
        RECT 51.900 168.040 53.100 168.340 ;
        RECT 54.890 168.070 56.000 168.340 ;
        RECT 60.120 168.070 60.620 174.110 ;
        RECT 63.860 174.100 65.420 174.110 ;
        RECT 64.360 173.870 65.420 174.100 ;
        RECT 67.640 173.970 69.140 174.570 ;
        RECT 71.530 174.100 77.160 174.600 ;
        RECT 83.070 174.410 84.870 174.710 ;
        RECT 87.570 174.410 89.370 174.710 ;
        RECT 83.070 174.110 84.270 174.410 ;
        RECT 88.170 174.110 89.370 174.410 ;
        RECT 67.040 173.670 68.240 173.970 ;
        RECT 68.540 173.670 69.740 173.970 ;
        RECT 71.530 173.870 72.640 174.100 ;
        RECT 83.070 173.810 83.970 174.110 ;
        RECT 88.470 173.810 89.370 174.110 ;
        RECT 65.540 173.370 67.640 173.670 ;
        RECT 69.140 173.370 71.540 173.670 ;
        RECT 83.370 173.510 83.670 173.810 ;
        RECT 85.170 173.510 85.470 173.810 ;
        RECT 85.770 173.510 86.070 173.810 ;
        RECT 86.370 173.510 86.670 173.810 ;
        RECT 86.970 173.510 87.270 173.810 ;
        RECT 88.770 173.510 89.070 173.810 ;
        RECT 65.240 173.070 67.040 173.370 ;
        RECT 69.740 173.070 71.540 173.370 ;
        RECT 65.240 172.770 66.440 173.070 ;
        RECT 70.340 172.770 71.540 173.070 ;
        RECT 85.170 172.910 87.270 173.510 ;
        RECT 65.240 172.470 66.140 172.770 ;
        RECT 70.640 172.470 71.540 172.770 ;
        RECT 84.870 172.610 85.770 172.910 ;
        RECT 86.670 172.610 87.870 172.910 ;
        RECT 65.540 172.170 65.840 172.470 ;
        RECT 67.340 172.170 67.640 172.470 ;
        RECT 67.940 172.170 68.240 172.470 ;
        RECT 68.540 172.170 68.840 172.470 ;
        RECT 69.140 172.170 69.440 172.470 ;
        RECT 70.940 172.170 71.240 172.470 ;
        RECT 84.270 172.310 86.070 172.610 ;
        RECT 86.370 172.310 87.870 172.610 ;
        RECT 67.340 171.570 69.440 172.170 ;
        RECT 84.270 172.010 84.870 172.310 ;
        RECT 85.470 172.010 86.970 172.310 ;
        RECT 87.570 172.010 88.170 172.310 ;
        RECT 84.270 171.710 84.570 172.010 ;
        RECT 67.040 171.270 67.940 171.570 ;
        RECT 68.840 171.270 70.040 171.570 ;
        RECT 66.440 170.970 68.240 171.270 ;
        RECT 68.540 170.970 70.040 171.270 ;
        RECT 83.970 171.410 84.570 171.710 ;
        RECT 83.970 171.110 84.870 171.410 ;
        RECT 85.770 171.110 86.670 172.010 ;
        RECT 87.870 171.710 88.170 172.010 ;
        RECT 94.590 171.960 95.090 175.440 ;
        RECT 101.710 175.230 102.010 175.530 ;
        RECT 103.210 175.230 104.110 176.130 ;
        RECT 105.010 175.830 105.910 176.130 ;
        RECT 105.310 175.530 105.910 175.830 ;
        RECT 105.310 175.230 105.610 175.530 ;
        RECT 101.710 174.930 102.310 175.230 ;
        RECT 102.910 174.930 104.410 175.230 ;
        RECT 105.010 174.930 105.610 175.230 ;
        RECT 101.710 174.630 103.510 174.930 ;
        RECT 103.810 174.630 105.310 174.930 ;
        RECT 102.310 174.330 103.210 174.630 ;
        RECT 104.110 174.330 105.310 174.630 ;
        RECT 102.610 173.730 104.710 174.330 ;
        RECT 100.810 173.430 101.710 173.730 ;
        RECT 102.610 173.430 102.910 173.730 ;
        RECT 103.210 173.430 103.510 173.730 ;
        RECT 103.810 173.430 104.110 173.730 ;
        RECT 104.410 173.430 104.710 173.730 ;
        RECT 105.610 173.430 106.510 173.730 ;
        RECT 100.510 172.830 102.010 173.430 ;
        RECT 105.310 172.830 106.810 173.430 ;
        RECT 100.810 172.530 102.610 172.830 ;
        RECT 104.710 172.530 106.510 172.830 ;
        RECT 101.710 172.230 102.910 172.530 ;
        RECT 104.410 172.230 105.610 172.530 ;
        RECT 99.630 171.960 100.690 172.230 ;
        RECT 87.870 171.410 88.470 171.710 ;
        RECT 94.590 171.460 100.690 171.960 ;
        RECT 102.310 171.930 103.510 172.230 ;
        RECT 103.810 171.930 105.010 172.230 ;
        RECT 106.800 171.960 107.910 172.230 ;
        RECT 87.570 171.110 88.470 171.410 ;
        RECT 99.630 171.230 100.690 171.460 ;
        RECT 102.910 171.330 104.410 171.930 ;
        RECT 106.800 171.460 111.190 171.960 ;
        RECT 66.440 170.670 67.040 170.970 ;
        RECT 67.640 170.670 69.140 170.970 ;
        RECT 69.740 170.670 70.340 170.970 ;
        RECT 66.440 170.370 66.740 170.670 ;
        RECT 66.140 170.070 66.740 170.370 ;
        RECT 66.140 169.770 67.040 170.070 ;
        RECT 67.940 169.770 68.840 170.670 ;
        RECT 70.040 170.370 70.340 170.670 ;
        RECT 70.040 170.070 70.640 170.370 ;
        RECT 69.740 169.770 70.640 170.070 ;
        RECT 83.970 169.910 88.470 171.110 ;
        RECT 102.310 171.030 103.510 171.330 ;
        RECT 103.810 171.030 105.010 171.330 ;
        RECT 106.800 171.230 107.910 171.460 ;
        RECT 100.810 170.730 102.910 171.030 ;
        RECT 104.410 170.730 106.810 171.030 ;
        RECT 100.510 170.430 102.310 170.730 ;
        RECT 105.010 170.430 106.810 170.730 ;
        RECT 100.510 170.130 101.710 170.430 ;
        RECT 105.610 170.130 106.810 170.430 ;
        RECT 66.140 168.570 70.640 169.770 ;
        RECT 82.690 169.270 84.080 169.710 ;
        RECT 84.270 169.310 88.170 169.910 ;
        RECT 100.510 169.830 101.410 170.130 ;
        RECT 105.910 169.830 106.810 170.130 ;
        RECT 100.810 169.530 101.110 169.830 ;
        RECT 102.610 169.530 102.910 169.830 ;
        RECT 103.210 169.530 103.510 169.830 ;
        RECT 103.810 169.530 104.110 169.830 ;
        RECT 104.410 169.530 104.710 169.830 ;
        RECT 106.210 169.530 106.510 169.830 ;
        RECT 82.690 169.100 83.250 169.270 ;
        RECT 84.870 169.010 87.570 169.310 ;
        RECT 85.170 168.710 87.570 169.010 ;
        RECT 102.610 168.930 104.710 169.530 ;
        RECT 102.310 168.630 103.210 168.930 ;
        RECT 104.110 168.630 105.310 168.930 ;
        RECT 36.710 163.190 39.110 163.490 ;
        RECT 34.230 162.920 34.680 163.030 ;
        RECT 34.230 162.420 35.340 162.920 ;
        RECT 36.410 162.890 39.110 163.190 ;
        RECT 35.810 162.290 39.710 162.890 ;
        RECT 35.510 161.090 40.010 162.290 ;
        RECT 35.510 160.790 36.410 161.090 ;
        RECT 35.510 160.490 36.110 160.790 ;
        RECT 35.810 160.190 36.110 160.490 ;
        RECT 37.310 160.190 38.210 161.090 ;
        RECT 39.110 160.790 40.010 161.090 ;
        RECT 39.410 160.490 40.010 160.790 ;
        RECT 39.410 160.190 39.710 160.490 ;
        RECT 35.810 159.890 36.410 160.190 ;
        RECT 37.010 159.890 38.510 160.190 ;
        RECT 39.110 159.890 39.710 160.190 ;
        RECT 35.810 159.590 37.610 159.890 ;
        RECT 37.910 159.590 39.410 159.890 ;
        RECT 36.410 159.290 37.310 159.590 ;
        RECT 38.210 159.290 39.410 159.590 ;
        RECT 36.710 158.690 38.810 159.290 ;
        RECT 34.910 158.390 35.810 158.690 ;
        RECT 36.710 158.390 37.010 158.690 ;
        RECT 37.310 158.390 37.610 158.690 ;
        RECT 37.910 158.390 38.210 158.690 ;
        RECT 38.510 158.390 38.810 158.690 ;
        RECT 39.710 158.390 40.610 158.690 ;
        RECT 34.610 157.790 36.110 158.390 ;
        RECT 39.410 157.790 40.910 158.390 ;
        RECT 34.910 157.490 36.710 157.790 ;
        RECT 38.810 157.490 40.610 157.790 ;
        RECT 35.810 157.190 37.010 157.490 ;
        RECT 38.510 157.190 39.710 157.490 ;
        RECT 33.730 156.920 34.790 157.190 ;
        RECT 31.830 156.420 34.790 156.920 ;
        RECT 36.410 156.890 37.610 157.190 ;
        RECT 37.910 156.890 39.110 157.190 ;
        RECT 40.900 156.920 42.010 157.190 ;
        RECT 44.210 156.920 44.710 167.590 ;
        RECT 47.220 167.570 48.780 167.590 ;
        RECT 47.720 167.340 48.780 167.570 ;
        RECT 51.000 167.440 52.500 168.040 ;
        RECT 54.890 167.570 60.620 168.070 ;
        RECT 64.860 167.930 66.250 168.370 ;
        RECT 66.440 167.970 70.340 168.570 ;
        RECT 101.710 168.330 103.510 168.630 ;
        RECT 103.810 168.330 105.310 168.630 ;
        RECT 101.710 168.030 102.310 168.330 ;
        RECT 102.910 168.030 104.410 168.330 ;
        RECT 105.010 168.030 105.610 168.330 ;
        RECT 64.860 167.760 65.420 167.930 ;
        RECT 67.040 167.670 69.740 167.970 ;
        RECT 101.710 167.730 102.010 168.030 ;
        RECT 50.400 167.140 51.600 167.440 ;
        RECT 51.900 167.140 53.100 167.440 ;
        RECT 54.890 167.340 56.000 167.570 ;
        RECT 67.340 167.370 69.740 167.670 ;
        RECT 101.410 167.430 102.010 167.730 ;
        RECT 48.900 166.840 51.000 167.140 ;
        RECT 52.500 166.840 54.900 167.140 ;
        RECT 48.600 166.540 50.400 166.840 ;
        RECT 53.100 166.540 54.900 166.840 ;
        RECT 48.600 166.240 49.800 166.540 ;
        RECT 53.700 166.240 54.900 166.540 ;
        RECT 48.600 165.940 49.500 166.240 ;
        RECT 54.000 165.940 54.900 166.240 ;
        RECT 101.410 167.130 102.310 167.430 ;
        RECT 103.210 167.130 104.110 168.030 ;
        RECT 105.310 167.730 105.610 168.030 ;
        RECT 105.310 167.430 105.910 167.730 ;
        RECT 105.010 167.130 105.910 167.430 ;
        RECT 48.900 165.640 49.200 165.940 ;
        RECT 50.700 165.640 51.000 165.940 ;
        RECT 51.300 165.640 51.600 165.940 ;
        RECT 51.900 165.640 52.200 165.940 ;
        RECT 52.500 165.640 52.800 165.940 ;
        RECT 54.300 165.640 54.600 165.940 ;
        RECT 101.410 165.930 105.910 167.130 ;
        RECT 50.700 165.040 52.800 165.640 ;
        RECT 100.130 165.290 101.520 165.730 ;
        RECT 101.710 165.330 105.610 165.930 ;
        RECT 100.130 165.120 100.690 165.290 ;
        RECT 50.400 164.740 51.300 165.040 ;
        RECT 52.200 164.740 53.400 165.040 ;
        RECT 102.310 165.030 105.010 165.330 ;
        RECT 49.800 164.440 51.600 164.740 ;
        RECT 51.900 164.440 53.400 164.740 ;
        RECT 102.610 164.730 105.010 165.030 ;
        RECT 49.800 164.140 50.400 164.440 ;
        RECT 51.000 164.140 52.500 164.440 ;
        RECT 53.100 164.140 53.700 164.440 ;
        RECT 49.800 163.840 50.100 164.140 ;
        RECT 49.500 163.540 50.100 163.840 ;
        RECT 49.500 163.240 50.400 163.540 ;
        RECT 51.300 163.240 52.200 164.140 ;
        RECT 53.400 163.840 53.700 164.140 ;
        RECT 53.400 163.540 54.000 163.840 ;
        RECT 53.100 163.240 54.000 163.540 ;
        RECT 49.500 162.040 54.000 163.240 ;
        RECT 110.690 163.010 111.190 171.460 ;
        RECT 118.090 169.280 120.490 169.580 ;
        RECT 115.610 169.010 116.060 169.120 ;
        RECT 115.610 168.510 116.720 169.010 ;
        RECT 117.790 168.980 120.490 169.280 ;
        RECT 117.190 168.380 121.090 168.980 ;
        RECT 116.890 167.180 121.390 168.380 ;
        RECT 116.890 166.880 117.790 167.180 ;
        RECT 116.890 166.580 117.490 166.880 ;
        RECT 117.190 166.280 117.490 166.580 ;
        RECT 118.690 166.280 119.590 167.180 ;
        RECT 120.490 166.880 121.390 167.180 ;
        RECT 120.790 166.580 121.390 166.880 ;
        RECT 120.790 166.280 121.090 166.580 ;
        RECT 117.190 165.980 117.790 166.280 ;
        RECT 118.390 165.980 119.890 166.280 ;
        RECT 120.490 165.980 121.090 166.280 ;
        RECT 117.190 165.680 118.990 165.980 ;
        RECT 119.290 165.680 120.790 165.980 ;
        RECT 117.790 165.380 118.690 165.680 ;
        RECT 119.590 165.380 120.790 165.680 ;
        RECT 118.090 164.780 120.190 165.380 ;
        RECT 116.290 164.480 117.190 164.780 ;
        RECT 118.090 164.480 118.390 164.780 ;
        RECT 118.690 164.480 118.990 164.780 ;
        RECT 119.290 164.480 119.590 164.780 ;
        RECT 119.890 164.480 120.190 164.780 ;
        RECT 121.090 164.480 121.990 164.780 ;
        RECT 115.990 163.880 117.490 164.480 ;
        RECT 120.790 163.880 122.290 164.480 ;
        RECT 116.290 163.580 118.090 163.880 ;
        RECT 120.190 163.580 121.990 163.880 ;
        RECT 117.190 163.280 118.390 163.580 ;
        RECT 119.890 163.280 121.090 163.580 ;
        RECT 115.110 163.010 116.170 163.280 ;
        RECT 110.690 162.510 116.170 163.010 ;
        RECT 117.790 162.980 118.990 163.280 ;
        RECT 119.290 162.980 120.490 163.280 ;
        RECT 122.280 163.020 123.390 163.280 ;
        RECT 115.110 162.280 116.170 162.510 ;
        RECT 118.390 162.380 119.890 162.980 ;
        RECT 122.280 162.520 127.280 163.020 ;
        RECT 122.280 162.510 123.780 162.520 ;
        RECT 117.790 162.080 118.990 162.380 ;
        RECT 119.290 162.080 120.490 162.380 ;
        RECT 122.280 162.280 123.390 162.510 ;
        RECT 48.220 161.400 49.610 161.840 ;
        RECT 49.800 161.440 53.700 162.040 ;
        RECT 116.290 161.780 118.390 162.080 ;
        RECT 119.890 161.780 122.290 162.080 ;
        RECT 115.990 161.480 117.790 161.780 ;
        RECT 120.490 161.480 122.290 161.780 ;
        RECT 48.220 161.230 48.780 161.400 ;
        RECT 50.400 161.140 53.100 161.440 ;
        RECT 50.700 160.840 53.100 161.140 ;
        RECT 115.990 161.180 117.190 161.480 ;
        RECT 121.090 161.180 122.290 161.480 ;
        RECT 115.990 160.880 116.890 161.180 ;
        RECT 121.390 160.880 122.290 161.180 ;
        RECT 116.290 160.580 116.590 160.880 ;
        RECT 118.090 160.580 118.390 160.880 ;
        RECT 118.690 160.580 118.990 160.880 ;
        RECT 119.290 160.580 119.590 160.880 ;
        RECT 119.890 160.580 120.190 160.880 ;
        RECT 121.690 160.580 121.990 160.880 ;
        RECT 118.090 159.980 120.190 160.580 ;
        RECT 117.790 159.680 118.690 159.980 ;
        RECT 119.590 159.680 120.790 159.980 ;
        RECT 117.190 159.380 118.990 159.680 ;
        RECT 119.290 159.380 120.790 159.680 ;
        RECT 117.190 159.080 117.790 159.380 ;
        RECT 118.390 159.080 119.890 159.380 ;
        RECT 120.490 159.080 121.090 159.380 ;
        RECT 117.190 158.780 117.490 159.080 ;
        RECT 116.890 158.480 117.490 158.780 ;
        RECT 116.890 158.180 117.790 158.480 ;
        RECT 118.690 158.180 119.590 159.080 ;
        RECT 120.790 158.780 121.090 159.080 ;
        RECT 120.790 158.480 121.390 158.780 ;
        RECT 120.490 158.180 121.390 158.480 ;
        RECT 116.890 156.980 121.390 158.180 ;
        RECT 26.640 148.410 29.040 148.710 ;
        RECT 24.160 148.140 24.610 148.250 ;
        RECT 24.160 147.640 25.270 148.140 ;
        RECT 26.340 148.110 29.040 148.410 ;
        RECT 25.740 147.510 29.640 148.110 ;
        RECT 25.440 146.310 29.940 147.510 ;
        RECT 25.440 146.010 26.340 146.310 ;
        RECT 25.440 145.710 26.040 146.010 ;
        RECT 25.740 145.410 26.040 145.710 ;
        RECT 27.240 145.410 28.140 146.310 ;
        RECT 29.040 146.010 29.940 146.310 ;
        RECT 29.340 145.710 29.940 146.010 ;
        RECT 29.340 145.410 29.640 145.710 ;
        RECT 25.740 145.110 26.340 145.410 ;
        RECT 26.940 145.110 28.440 145.410 ;
        RECT 29.040 145.110 29.640 145.410 ;
        RECT 25.740 144.810 27.540 145.110 ;
        RECT 27.840 144.810 29.340 145.110 ;
        RECT 26.340 144.510 27.240 144.810 ;
        RECT 28.140 144.510 29.340 144.810 ;
        RECT 26.640 143.910 28.740 144.510 ;
        RECT 24.840 143.610 25.740 143.910 ;
        RECT 26.640 143.610 26.940 143.910 ;
        RECT 27.240 143.610 27.540 143.910 ;
        RECT 27.840 143.610 28.140 143.910 ;
        RECT 28.440 143.610 28.740 143.910 ;
        RECT 29.640 143.610 30.540 143.910 ;
        RECT 24.540 143.010 26.040 143.610 ;
        RECT 29.340 143.010 30.840 143.610 ;
        RECT 24.840 142.710 26.640 143.010 ;
        RECT 28.740 142.710 30.540 143.010 ;
        RECT 25.740 142.410 26.940 142.710 ;
        RECT 28.440 142.410 29.640 142.710 ;
        RECT 31.830 142.410 32.330 156.420 ;
        RECT 33.730 156.190 34.790 156.420 ;
        RECT 37.010 156.290 38.510 156.890 ;
        RECT 40.900 156.420 44.710 156.920 ;
        RECT 36.410 155.990 37.610 156.290 ;
        RECT 37.910 155.990 39.110 156.290 ;
        RECT 40.900 156.190 42.010 156.420 ;
        RECT 115.610 156.340 117.000 156.780 ;
        RECT 117.190 156.380 121.090 156.980 ;
        RECT 115.610 156.170 116.170 156.340 ;
        RECT 117.790 156.080 120.490 156.380 ;
        RECT 34.910 155.690 37.010 155.990 ;
        RECT 38.510 155.690 40.910 155.990 ;
        RECT 118.090 155.780 120.490 156.080 ;
        RECT 34.610 155.390 36.410 155.690 ;
        RECT 39.110 155.390 40.910 155.690 ;
        RECT 34.610 155.090 35.810 155.390 ;
        RECT 39.710 155.090 40.910 155.390 ;
        RECT 34.610 154.790 35.510 155.090 ;
        RECT 40.010 154.790 40.910 155.090 ;
        RECT 34.910 154.490 35.210 154.790 ;
        RECT 36.710 154.490 37.010 154.790 ;
        RECT 37.310 154.490 37.610 154.790 ;
        RECT 37.910 154.490 38.210 154.790 ;
        RECT 38.510 154.490 38.810 154.790 ;
        RECT 40.310 154.490 40.610 154.790 ;
        RECT 36.710 153.890 38.810 154.490 ;
        RECT 36.410 153.590 37.310 153.890 ;
        RECT 38.210 153.590 39.410 153.890 ;
        RECT 35.810 153.290 37.610 153.590 ;
        RECT 37.910 153.290 39.410 153.590 ;
        RECT 35.810 152.990 36.410 153.290 ;
        RECT 37.010 152.990 38.510 153.290 ;
        RECT 39.110 152.990 39.710 153.290 ;
        RECT 35.810 152.690 36.110 152.990 ;
        RECT 35.510 152.390 36.110 152.690 ;
        RECT 35.510 152.090 36.410 152.390 ;
        RECT 37.310 152.090 38.210 152.990 ;
        RECT 39.410 152.690 39.710 152.990 ;
        RECT 39.410 152.390 40.010 152.690 ;
        RECT 39.110 152.090 40.010 152.390 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 35.510 150.890 40.010 152.090 ;
        RECT 34.230 150.250 35.620 150.690 ;
        RECT 35.810 150.290 39.710 150.890 ;
        RECT 34.230 150.080 34.790 150.250 ;
        RECT 36.410 149.990 39.110 150.290 ;
        RECT 36.710 149.690 39.110 149.990 ;
        RECT 68.170 149.600 91.570 152.200 ;
        RECT 126.780 150.170 127.280 162.520 ;
        RECT 130.260 156.170 132.660 156.470 ;
        RECT 127.780 155.900 128.230 156.010 ;
        RECT 127.780 155.400 128.890 155.900 ;
        RECT 129.960 155.870 132.660 156.170 ;
        RECT 129.360 155.270 133.260 155.870 ;
        RECT 129.060 154.070 133.560 155.270 ;
        RECT 129.060 153.770 129.960 154.070 ;
        RECT 129.060 153.470 129.660 153.770 ;
        RECT 129.360 153.170 129.660 153.470 ;
        RECT 130.860 153.170 131.760 154.070 ;
        RECT 132.660 153.770 133.560 154.070 ;
        RECT 132.960 153.470 133.560 153.770 ;
        RECT 132.960 153.170 133.260 153.470 ;
        RECT 129.360 152.870 129.960 153.170 ;
        RECT 130.560 152.870 132.060 153.170 ;
        RECT 132.660 152.870 133.260 153.170 ;
        RECT 129.360 152.570 131.160 152.870 ;
        RECT 131.460 152.570 132.960 152.870 ;
        RECT 129.960 152.270 130.860 152.570 ;
        RECT 131.760 152.270 132.960 152.570 ;
        RECT 130.260 151.670 132.360 152.270 ;
        RECT 128.460 151.370 129.360 151.670 ;
        RECT 130.260 151.370 130.560 151.670 ;
        RECT 130.860 151.370 131.160 151.670 ;
        RECT 131.460 151.370 131.760 151.670 ;
        RECT 132.060 151.370 132.360 151.670 ;
        RECT 133.260 151.370 134.160 151.670 ;
        RECT 128.160 150.770 129.660 151.370 ;
        RECT 132.960 150.770 134.460 151.370 ;
        RECT 128.460 150.470 130.260 150.770 ;
        RECT 132.360 150.470 134.160 150.770 ;
        RECT 129.360 150.170 130.560 150.470 ;
        RECT 132.060 150.170 133.260 150.470 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 126.780 149.400 128.340 150.170 ;
        RECT 129.960 149.870 131.160 150.170 ;
        RECT 131.460 149.870 132.660 150.170 ;
        RECT 134.450 149.900 135.560 150.170 ;
        RECT 127.280 149.170 128.340 149.400 ;
        RECT 130.560 149.270 132.060 149.870 ;
        RECT 134.450 149.850 135.950 149.900 ;
        RECT 129.960 148.970 131.160 149.270 ;
        RECT 131.460 148.970 132.660 149.270 ;
        RECT 134.450 149.170 135.970 149.850 ;
        RECT 128.460 148.670 130.560 148.970 ;
        RECT 132.060 148.670 134.460 148.970 ;
        RECT 128.160 148.370 129.960 148.670 ;
        RECT 132.660 148.370 134.460 148.670 ;
        RECT 128.160 148.070 129.360 148.370 ;
        RECT 133.260 148.070 134.460 148.370 ;
        RECT 128.160 147.770 129.060 148.070 ;
        RECT 133.560 147.770 134.460 148.070 ;
        RECT 128.460 147.470 128.760 147.770 ;
        RECT 130.260 147.470 130.560 147.770 ;
        RECT 130.860 147.470 131.160 147.770 ;
        RECT 131.460 147.470 131.760 147.770 ;
        RECT 132.060 147.470 132.360 147.770 ;
        RECT 133.860 147.470 134.160 147.770 ;
        RECT 130.260 146.870 132.360 147.470 ;
        RECT 129.960 146.570 130.860 146.870 ;
        RECT 131.760 146.570 132.960 146.870 ;
        RECT 129.360 146.270 131.160 146.570 ;
        RECT 131.460 146.270 132.960 146.570 ;
        RECT 129.360 145.970 129.960 146.270 ;
        RECT 130.560 145.970 132.060 146.270 ;
        RECT 132.660 145.970 133.260 146.270 ;
        RECT 129.360 145.670 129.660 145.970 ;
        RECT 129.060 145.370 129.660 145.670 ;
        RECT 129.060 145.070 129.960 145.370 ;
        RECT 130.860 145.070 131.760 145.970 ;
        RECT 132.960 145.670 133.260 145.970 ;
        RECT 135.470 146.060 135.970 149.170 ;
        RECT 132.960 145.370 133.560 145.670 ;
        RECT 135.470 145.560 141.000 146.060 ;
        RECT 132.660 145.070 133.560 145.370 ;
        RECT 23.660 142.140 24.720 142.410 ;
        RECT 23.160 141.410 24.720 142.140 ;
        RECT 26.340 142.110 27.540 142.410 ;
        RECT 27.840 142.110 29.040 142.410 ;
        RECT 26.940 141.510 28.440 142.110 ;
        RECT 30.830 141.640 32.330 142.410 ;
        RECT 23.160 134.340 23.660 141.410 ;
        RECT 26.340 141.210 27.540 141.510 ;
        RECT 27.840 141.210 29.040 141.510 ;
        RECT 30.830 141.410 31.940 141.640 ;
        RECT 24.840 140.910 26.940 141.210 ;
        RECT 28.440 140.910 30.840 141.210 ;
        RECT 24.540 140.610 26.340 140.910 ;
        RECT 29.040 140.610 30.840 140.910 ;
        RECT 24.540 140.310 25.740 140.610 ;
        RECT 29.640 140.310 30.840 140.610 ;
        RECT 24.540 140.010 25.440 140.310 ;
        RECT 29.940 140.010 30.840 140.310 ;
        RECT 24.840 139.710 25.140 140.010 ;
        RECT 26.640 139.710 26.940 140.010 ;
        RECT 27.240 139.710 27.540 140.010 ;
        RECT 27.840 139.710 28.140 140.010 ;
        RECT 28.440 139.710 28.740 140.010 ;
        RECT 30.240 139.710 30.540 140.010 ;
        RECT 26.640 139.110 28.740 139.710 ;
        RECT 26.340 138.810 27.240 139.110 ;
        RECT 28.140 138.810 29.340 139.110 ;
        RECT 25.740 138.510 27.540 138.810 ;
        RECT 27.840 138.510 29.340 138.810 ;
        RECT 25.740 138.210 26.340 138.510 ;
        RECT 26.940 138.210 28.440 138.510 ;
        RECT 29.040 138.210 29.640 138.510 ;
        RECT 25.740 137.910 26.040 138.210 ;
        RECT 25.440 137.610 26.040 137.910 ;
        RECT 25.440 137.310 26.340 137.610 ;
        RECT 27.240 137.310 28.140 138.210 ;
        RECT 29.340 137.910 29.640 138.210 ;
        RECT 29.340 137.610 29.940 137.910 ;
        RECT 29.040 137.310 29.940 137.610 ;
        RECT 25.440 136.110 29.940 137.310 ;
        RECT 24.160 135.470 25.550 135.910 ;
        RECT 25.740 135.510 29.640 136.110 ;
        RECT 24.160 135.300 24.720 135.470 ;
        RECT 26.340 135.210 29.040 135.510 ;
        RECT 26.640 134.910 29.040 135.210 ;
        RECT 15.180 133.840 23.660 134.340 ;
        RECT 60.370 134.000 99.370 144.400 ;
        RECT 129.060 143.870 133.560 145.070 ;
        RECT 127.780 143.230 129.170 143.670 ;
        RECT 129.360 143.270 133.260 143.870 ;
        RECT 127.780 143.060 128.340 143.230 ;
        RECT 129.960 142.970 132.660 143.270 ;
        RECT 130.260 142.670 132.660 142.970 ;
        RECT 135.120 140.060 137.520 140.360 ;
        RECT 135.120 139.760 137.820 140.060 ;
        RECT 139.550 139.790 140.000 139.900 ;
        RECT 134.520 139.160 138.420 139.760 ;
        RECT 138.890 139.290 140.000 139.790 ;
        RECT 134.220 137.960 138.720 139.160 ;
        RECT 134.220 137.660 135.120 137.960 ;
        RECT 134.220 137.360 134.820 137.660 ;
        RECT 134.520 137.060 134.820 137.360 ;
        RECT 136.020 137.060 136.920 137.960 ;
        RECT 137.820 137.660 138.720 137.960 ;
        RECT 138.120 137.360 138.720 137.660 ;
        RECT 138.120 137.060 138.420 137.360 ;
        RECT 134.520 136.760 135.120 137.060 ;
        RECT 135.720 136.760 137.220 137.060 ;
        RECT 137.820 136.760 138.420 137.060 ;
        RECT 134.820 136.460 136.320 136.760 ;
        RECT 136.620 136.460 138.420 136.760 ;
        RECT 134.820 136.160 136.020 136.460 ;
        RECT 136.920 136.160 137.820 136.460 ;
        RECT 135.420 135.560 137.520 136.160 ;
        RECT 133.620 135.260 134.520 135.560 ;
        RECT 135.420 135.260 135.720 135.560 ;
        RECT 136.020 135.260 136.320 135.560 ;
        RECT 136.620 135.260 136.920 135.560 ;
        RECT 137.220 135.260 137.520 135.560 ;
        RECT 138.420 135.260 139.320 135.560 ;
        RECT 133.320 134.660 134.820 135.260 ;
        RECT 138.120 134.660 139.620 135.260 ;
        RECT 133.620 134.360 135.420 134.660 ;
        RECT 137.520 134.360 139.320 134.660 ;
        RECT 134.520 134.060 135.720 134.360 ;
        RECT 137.220 134.060 138.420 134.360 ;
        RECT 140.500 134.060 141.000 145.560 ;
        RECT 15.180 125.320 15.680 133.840 ;
        RECT 18.470 131.320 20.870 131.620 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 18.470 131.020 21.170 131.320 ;
        RECT 22.900 131.050 23.350 131.160 ;
        RECT 17.870 130.420 21.770 131.020 ;
        RECT 22.240 130.550 23.350 131.050 ;
        RECT 17.570 129.220 22.070 130.420 ;
        RECT 17.570 128.920 18.470 129.220 ;
        RECT 17.570 128.620 18.170 128.920 ;
        RECT 17.870 128.320 18.170 128.620 ;
        RECT 19.370 128.320 20.270 129.220 ;
        RECT 21.170 128.920 22.070 129.220 ;
        RECT 21.470 128.620 22.070 128.920 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 21.470 128.320 21.770 128.620 ;
        RECT 17.870 128.020 18.470 128.320 ;
        RECT 19.070 128.020 20.570 128.320 ;
        RECT 21.170 128.020 21.770 128.320 ;
        RECT 18.170 127.720 19.670 128.020 ;
        RECT 19.970 127.720 21.770 128.020 ;
        RECT 18.170 127.420 19.370 127.720 ;
        RECT 20.270 127.420 21.170 127.720 ;
        RECT 18.770 126.820 20.870 127.420 ;
        RECT 16.970 126.520 17.870 126.820 ;
        RECT 18.770 126.520 19.070 126.820 ;
        RECT 19.370 126.520 19.670 126.820 ;
        RECT 19.970 126.520 20.270 126.820 ;
        RECT 20.570 126.520 20.870 126.820 ;
        RECT 21.770 126.520 22.670 126.820 ;
        RECT 16.670 125.920 18.170 126.520 ;
        RECT 21.470 125.920 22.970 126.520 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 132.220 133.790 133.330 134.060 ;
        RECT 131.830 133.750 133.330 133.790 ;
        RECT 135.120 133.760 136.320 134.060 ;
        RECT 136.620 133.760 137.820 134.060 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 131.820 133.060 133.330 133.750 ;
        RECT 135.720 133.160 137.220 133.760 ;
        RECT 139.440 133.290 141.000 134.060 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 16.970 125.620 18.770 125.920 ;
        RECT 20.870 125.620 22.670 125.920 ;
        RECT 17.870 125.320 19.070 125.620 ;
        RECT 20.570 125.320 21.770 125.620 ;
        RECT 15.180 124.550 16.680 125.320 ;
        RECT 18.470 125.020 19.670 125.320 ;
        RECT 19.970 125.020 21.170 125.320 ;
        RECT 22.790 125.050 23.850 125.320 ;
        RECT 22.790 125.040 24.350 125.050 ;
        RECT 15.570 124.320 16.680 124.550 ;
        RECT 19.070 124.420 20.570 125.020 ;
        RECT 22.790 124.540 27.060 125.040 ;
        RECT 18.470 124.120 19.670 124.420 ;
        RECT 19.970 124.120 21.170 124.420 ;
        RECT 22.790 124.320 23.850 124.540 ;
        RECT 16.670 123.820 19.070 124.120 ;
        RECT 20.570 123.820 22.670 124.120 ;
        RECT 16.670 123.520 18.470 123.820 ;
        RECT 21.170 123.520 22.970 123.820 ;
        RECT 16.670 123.220 17.870 123.520 ;
        RECT 21.770 123.220 22.970 123.520 ;
        RECT 16.670 122.920 17.570 123.220 ;
        RECT 22.070 122.920 22.970 123.220 ;
        RECT 16.970 122.620 17.270 122.920 ;
        RECT 18.770 122.620 19.070 122.920 ;
        RECT 19.370 122.620 19.670 122.920 ;
        RECT 19.970 122.620 20.270 122.920 ;
        RECT 20.570 122.620 20.870 122.920 ;
        RECT 22.370 122.620 22.670 122.920 ;
        RECT 18.770 122.020 20.870 122.620 ;
        RECT 18.170 121.720 19.370 122.020 ;
        RECT 20.270 121.720 21.170 122.020 ;
        RECT 18.170 121.420 19.670 121.720 ;
        RECT 19.970 121.420 21.770 121.720 ;
        RECT 17.870 121.120 18.470 121.420 ;
        RECT 19.070 121.120 20.570 121.420 ;
        RECT 21.170 121.120 21.770 121.420 ;
        RECT 17.870 120.820 18.170 121.120 ;
        RECT 17.570 120.520 18.170 120.820 ;
        RECT 17.570 120.220 18.470 120.520 ;
        RECT 19.370 120.220 20.270 121.120 ;
        RECT 21.470 120.820 21.770 121.120 ;
        RECT 21.470 120.520 22.070 120.820 ;
        RECT 21.170 120.220 22.070 120.520 ;
        RECT 17.570 119.020 22.070 120.220 ;
        RECT 17.870 118.420 21.770 119.020 ;
        RECT 18.470 118.120 21.170 118.420 ;
        RECT 21.960 118.380 23.350 118.820 ;
        RECT 22.790 118.210 23.350 118.380 ;
        RECT 18.470 117.820 20.870 118.120 ;
        RECT 7.470 112.910 9.070 114.410 ;
        RECT 21.370 113.440 23.770 113.740 ;
        RECT 18.890 113.170 19.340 113.280 ;
        RECT 18.890 112.670 20.000 113.170 ;
        RECT 21.070 113.140 23.770 113.440 ;
        RECT 20.470 112.540 24.370 113.140 ;
        RECT 20.170 111.340 24.670 112.540 ;
        RECT 20.170 111.040 21.070 111.340 ;
        RECT 20.170 110.740 20.770 111.040 ;
        RECT 20.470 110.440 20.770 110.740 ;
        RECT 21.970 110.440 22.870 111.340 ;
        RECT 23.770 111.040 24.670 111.340 ;
        RECT 24.070 110.740 24.670 111.040 ;
        RECT 24.070 110.440 24.370 110.740 ;
        RECT 20.470 110.140 21.070 110.440 ;
        RECT 21.670 110.140 23.170 110.440 ;
        RECT 23.770 110.140 24.370 110.440 ;
        RECT 20.470 109.840 22.270 110.140 ;
        RECT 22.570 109.840 24.070 110.140 ;
        RECT 21.070 109.540 21.970 109.840 ;
        RECT 22.870 109.540 24.070 109.840 ;
        RECT 21.370 108.940 23.470 109.540 ;
        RECT 19.570 108.640 20.470 108.940 ;
        RECT 21.370 108.640 21.670 108.940 ;
        RECT 21.970 108.640 22.270 108.940 ;
        RECT 22.570 108.640 22.870 108.940 ;
        RECT 23.170 108.640 23.470 108.940 ;
        RECT 24.370 108.640 25.270 108.940 ;
        RECT 19.270 108.040 20.770 108.640 ;
        RECT 24.070 108.040 25.570 108.640 ;
        RECT 19.570 107.740 21.370 108.040 ;
        RECT 23.470 107.740 25.270 108.040 ;
        RECT 20.470 107.440 21.670 107.740 ;
        RECT 23.170 107.440 24.370 107.740 ;
        RECT 26.560 107.440 27.060 124.540 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 30.710 114.330 31.810 115.530 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 131.820 116.110 132.320 133.060 ;
        RECT 135.120 132.860 136.320 133.160 ;
        RECT 136.620 132.860 137.820 133.160 ;
        RECT 139.440 133.060 140.500 133.290 ;
        RECT 133.320 132.560 135.720 132.860 ;
        RECT 137.220 132.560 139.320 132.860 ;
        RECT 133.320 132.260 135.120 132.560 ;
        RECT 137.820 132.260 139.620 132.560 ;
        RECT 133.320 131.960 134.520 132.260 ;
        RECT 138.420 131.960 139.620 132.260 ;
        RECT 133.320 131.660 134.220 131.960 ;
        RECT 138.720 131.660 139.620 131.960 ;
        RECT 133.620 131.360 133.920 131.660 ;
        RECT 135.420 131.360 135.720 131.660 ;
        RECT 136.020 131.360 136.320 131.660 ;
        RECT 136.620 131.360 136.920 131.660 ;
        RECT 137.220 131.360 137.520 131.660 ;
        RECT 139.020 131.360 139.320 131.660 ;
        RECT 135.420 130.760 137.520 131.360 ;
        RECT 134.820 130.460 136.020 130.760 ;
        RECT 136.920 130.460 137.820 130.760 ;
        RECT 134.820 130.160 136.320 130.460 ;
        RECT 136.620 130.160 138.420 130.460 ;
        RECT 134.520 129.860 135.120 130.160 ;
        RECT 135.720 129.860 137.220 130.160 ;
        RECT 137.820 129.860 138.420 130.160 ;
        RECT 134.520 129.560 134.820 129.860 ;
        RECT 134.220 129.260 134.820 129.560 ;
        RECT 134.220 128.960 135.120 129.260 ;
        RECT 136.020 128.960 136.920 129.860 ;
        RECT 138.120 129.560 138.420 129.860 ;
        RECT 138.120 129.260 138.720 129.560 ;
        RECT 137.820 128.960 138.720 129.260 ;
        RECT 134.220 127.760 138.720 128.960 ;
        RECT 134.520 127.160 138.420 127.760 ;
        RECT 135.120 126.860 137.820 127.160 ;
        RECT 138.610 127.120 140.000 127.560 ;
        RECT 139.440 126.950 140.000 127.120 ;
        RECT 135.120 126.560 137.520 126.860 ;
        RECT 140.690 122.380 143.090 122.680 ;
        RECT 138.210 122.110 138.660 122.220 ;
        RECT 138.210 121.610 139.320 122.110 ;
        RECT 140.390 122.080 143.090 122.380 ;
        RECT 139.790 121.480 143.690 122.080 ;
        RECT 139.490 120.280 143.990 121.480 ;
        RECT 139.490 119.980 140.390 120.280 ;
        RECT 139.490 119.680 140.090 119.980 ;
        RECT 139.790 119.380 140.090 119.680 ;
        RECT 141.290 119.380 142.190 120.280 ;
        RECT 143.090 119.980 143.990 120.280 ;
        RECT 143.390 119.680 143.990 119.980 ;
        RECT 143.390 119.380 143.690 119.680 ;
        RECT 139.790 119.080 140.390 119.380 ;
        RECT 140.990 119.080 142.490 119.380 ;
        RECT 143.090 119.080 143.690 119.380 ;
        RECT 139.790 118.780 141.590 119.080 ;
        RECT 141.890 118.780 143.390 119.080 ;
        RECT 140.390 118.480 141.290 118.780 ;
        RECT 142.190 118.480 143.390 118.780 ;
        RECT 140.690 117.880 142.790 118.480 ;
        RECT 138.890 117.580 139.790 117.880 ;
        RECT 140.690 117.580 140.990 117.880 ;
        RECT 141.290 117.580 141.590 117.880 ;
        RECT 141.890 117.580 142.190 117.880 ;
        RECT 142.490 117.580 142.790 117.880 ;
        RECT 143.690 117.580 144.590 117.880 ;
        RECT 138.590 116.980 140.090 117.580 ;
        RECT 143.390 116.980 144.890 117.580 ;
        RECT 138.890 116.680 140.690 116.980 ;
        RECT 142.790 116.680 144.590 116.980 ;
        RECT 139.790 116.380 140.990 116.680 ;
        RECT 142.490 116.380 143.690 116.680 ;
        RECT 137.710 116.110 138.770 116.380 ;
        RECT 131.820 115.610 138.770 116.110 ;
        RECT 140.390 116.080 141.590 116.380 ;
        RECT 141.890 116.080 143.090 116.380 ;
        RECT 144.880 116.110 145.990 116.380 ;
        RECT 137.710 115.380 138.770 115.610 ;
        RECT 140.990 115.480 142.490 116.080 ;
        RECT 144.880 116.010 146.380 116.110 ;
        RECT 140.390 115.180 141.590 115.480 ;
        RECT 141.890 115.180 143.090 115.480 ;
        RECT 144.880 115.380 146.390 116.010 ;
        RECT 138.890 114.880 140.990 115.180 ;
        RECT 142.490 114.880 144.890 115.180 ;
        RECT 138.590 114.580 140.390 114.880 ;
        RECT 143.090 114.580 144.890 114.880 ;
        RECT 138.590 114.280 139.790 114.580 ;
        RECT 143.690 114.280 144.890 114.580 ;
        RECT 138.590 113.980 139.490 114.280 ;
        RECT 143.990 113.980 144.890 114.280 ;
        RECT 138.890 113.680 139.190 113.980 ;
        RECT 140.690 113.680 140.990 113.980 ;
        RECT 141.290 113.680 141.590 113.980 ;
        RECT 141.890 113.680 142.190 113.980 ;
        RECT 142.490 113.680 142.790 113.980 ;
        RECT 144.290 113.680 144.590 113.980 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 140.690 113.080 142.790 113.680 ;
        RECT 140.390 112.780 141.290 113.080 ;
        RECT 142.190 112.780 143.390 113.080 ;
        RECT 139.790 112.480 141.590 112.780 ;
        RECT 141.890 112.480 143.390 112.780 ;
        RECT 139.790 112.180 140.390 112.480 ;
        RECT 140.990 112.180 142.490 112.480 ;
        RECT 143.090 112.180 143.690 112.480 ;
        RECT 139.790 111.880 140.090 112.180 ;
        RECT 139.490 111.580 140.090 111.880 ;
        RECT 139.490 111.280 140.390 111.580 ;
        RECT 141.290 111.280 142.190 112.180 ;
        RECT 143.390 111.880 143.690 112.180 ;
        RECT 143.390 111.580 143.990 111.880 ;
        RECT 143.090 111.280 143.990 111.580 ;
        RECT 18.390 107.170 19.450 107.440 ;
        RECT 17.890 106.440 19.450 107.170 ;
        RECT 21.070 107.140 22.270 107.440 ;
        RECT 22.570 107.140 23.770 107.440 ;
        RECT 21.670 106.540 23.170 107.140 ;
        RECT 25.560 106.670 27.060 107.440 ;
        RECT 17.890 90.060 18.390 106.440 ;
        RECT 21.070 106.240 22.270 106.540 ;
        RECT 22.570 106.240 23.770 106.540 ;
        RECT 25.560 106.440 26.670 106.670 ;
        RECT 19.570 105.940 21.670 106.240 ;
        RECT 23.170 105.940 25.570 106.240 ;
        RECT 19.270 105.640 21.070 105.940 ;
        RECT 23.770 105.640 25.570 105.940 ;
        RECT 19.270 105.340 20.470 105.640 ;
        RECT 24.370 105.340 25.570 105.640 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
        RECT 139.490 110.080 143.990 111.280 ;
        RECT 138.210 109.440 139.600 109.880 ;
        RECT 139.790 109.480 143.690 110.080 ;
        RECT 138.210 109.270 138.770 109.440 ;
        RECT 140.390 109.180 143.090 109.480 ;
        RECT 140.690 108.880 143.090 109.180 ;
        RECT 19.270 105.040 20.170 105.340 ;
        RECT 24.670 105.040 25.570 105.340 ;
        RECT 19.570 104.740 19.870 105.040 ;
        RECT 21.370 104.740 21.670 105.040 ;
        RECT 21.970 104.740 22.270 105.040 ;
        RECT 22.570 104.740 22.870 105.040 ;
        RECT 23.170 104.740 23.470 105.040 ;
        RECT 24.970 104.740 25.270 105.040 ;
        RECT 21.370 104.140 23.470 104.740 ;
        RECT 21.070 103.840 21.970 104.140 ;
        RECT 22.870 103.840 24.070 104.140 ;
        RECT 20.470 103.540 22.270 103.840 ;
        RECT 22.570 103.540 24.070 103.840 ;
        RECT 20.470 103.240 21.070 103.540 ;
        RECT 21.670 103.240 23.170 103.540 ;
        RECT 23.770 103.240 24.370 103.540 ;
        RECT 20.470 102.940 20.770 103.240 ;
        RECT 20.170 102.640 20.770 102.940 ;
        RECT 20.170 102.340 21.070 102.640 ;
        RECT 21.970 102.340 22.870 103.240 ;
        RECT 24.070 102.940 24.370 103.240 ;
        RECT 24.070 102.640 24.670 102.940 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 135.120 104.700 137.520 105.000 ;
        RECT 135.120 104.400 137.820 104.700 ;
        RECT 139.550 104.430 140.000 104.540 ;
        RECT 134.520 103.800 138.420 104.400 ;
        RECT 138.890 103.930 140.000 104.430 ;
        RECT 23.770 102.340 24.670 102.640 ;
        RECT 20.170 101.140 24.670 102.340 ;
        RECT 18.890 100.500 20.280 100.940 ;
        RECT 20.470 100.540 24.370 101.140 ;
        RECT 18.890 100.330 19.450 100.500 ;
        RECT 21.070 100.240 23.770 100.540 ;
        RECT 21.370 99.940 23.770 100.240 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 134.220 102.600 138.720 103.800 ;
        RECT 134.220 102.300 135.120 102.600 ;
        RECT 134.220 102.000 134.820 102.300 ;
        RECT 134.520 101.700 134.820 102.000 ;
        RECT 136.020 101.700 136.920 102.600 ;
        RECT 137.820 102.300 138.720 102.600 ;
        RECT 138.120 102.000 138.720 102.300 ;
        RECT 138.120 101.700 138.420 102.000 ;
        RECT 134.520 101.400 135.120 101.700 ;
        RECT 135.720 101.400 137.220 101.700 ;
        RECT 137.820 101.400 138.420 101.700 ;
        RECT 134.820 101.100 136.320 101.400 ;
        RECT 136.620 101.100 138.420 101.400 ;
        RECT 134.820 100.800 136.020 101.100 ;
        RECT 136.920 100.800 137.820 101.100 ;
        RECT 135.420 100.200 137.520 100.800 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
        RECT 133.620 99.900 134.520 100.200 ;
        RECT 135.420 99.900 135.720 100.200 ;
        RECT 136.020 99.900 136.320 100.200 ;
        RECT 136.620 99.900 136.920 100.200 ;
        RECT 137.220 99.900 137.520 100.200 ;
        RECT 138.420 99.900 139.320 100.200 ;
        RECT 133.320 99.300 134.820 99.900 ;
        RECT 138.120 99.300 139.620 99.900 ;
        RECT 133.620 99.000 135.420 99.300 ;
        RECT 137.520 99.000 139.320 99.300 ;
        RECT 134.520 98.700 135.720 99.000 ;
        RECT 137.220 98.700 138.420 99.000 ;
        RECT 132.220 98.430 133.330 98.700 ;
        RECT 131.830 97.700 133.330 98.430 ;
        RECT 135.120 98.400 136.320 98.700 ;
        RECT 136.620 98.400 137.820 98.700 ;
        RECT 139.440 98.430 140.500 98.700 ;
        RECT 145.890 98.430 146.390 115.380 ;
        RECT 135.720 97.800 137.220 98.400 ;
        RECT 139.440 97.930 146.390 98.430 ;
        RECT 23.740 96.350 26.140 96.650 ;
        RECT 23.740 96.050 26.440 96.350 ;
        RECT 28.170 96.080 28.620 96.190 ;
        RECT 23.140 95.450 27.040 96.050 ;
        RECT 27.510 95.580 28.620 96.080 ;
        RECT 22.840 94.250 27.340 95.450 ;
        RECT 22.840 93.950 23.740 94.250 ;
        RECT 22.840 93.650 23.440 93.950 ;
        RECT 23.140 93.350 23.440 93.650 ;
        RECT 24.640 93.350 25.540 94.250 ;
        RECT 26.440 93.950 27.340 94.250 ;
        RECT 26.740 93.650 27.340 93.950 ;
        RECT 26.740 93.350 27.040 93.650 ;
        RECT 23.140 93.050 23.740 93.350 ;
        RECT 24.340 93.050 25.840 93.350 ;
        RECT 26.440 93.050 27.040 93.350 ;
        RECT 23.440 92.750 24.940 93.050 ;
        RECT 25.240 92.750 27.040 93.050 ;
        RECT 23.440 92.450 24.640 92.750 ;
        RECT 25.540 92.450 26.440 92.750 ;
        RECT 24.040 91.850 26.140 92.450 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 22.240 91.550 23.140 91.850 ;
        RECT 24.040 91.550 24.340 91.850 ;
        RECT 24.640 91.550 24.940 91.850 ;
        RECT 25.240 91.550 25.540 91.850 ;
        RECT 25.840 91.550 26.140 91.850 ;
        RECT 27.040 91.550 27.940 91.850 ;
        RECT 21.940 90.950 23.440 91.550 ;
        RECT 26.740 90.950 28.240 91.550 ;
        RECT 22.240 90.650 24.040 90.950 ;
        RECT 26.140 90.650 27.940 90.950 ;
        RECT 23.140 90.350 24.340 90.650 ;
        RECT 25.840 90.350 27.040 90.650 ;
        RECT 20.840 90.080 21.950 90.350 ;
        RECT 20.450 90.060 21.950 90.080 ;
        RECT 17.890 89.580 21.950 90.060 ;
        RECT 23.740 90.050 24.940 90.350 ;
        RECT 25.240 90.050 26.440 90.350 ;
        RECT 28.060 90.080 29.120 90.350 ;
        RECT 28.060 90.060 29.620 90.080 ;
        RECT 17.890 89.560 20.650 89.580 ;
        RECT 20.840 89.350 21.950 89.580 ;
        RECT 24.340 89.450 25.840 90.050 ;
        RECT 28.060 89.560 31.020 90.060 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
        RECT 131.830 90.060 132.330 97.700 ;
        RECT 135.120 97.500 136.320 97.800 ;
        RECT 136.620 97.500 137.820 97.800 ;
        RECT 139.440 97.700 140.500 97.930 ;
        RECT 133.320 97.200 135.720 97.500 ;
        RECT 137.220 97.200 139.320 97.500 ;
        RECT 133.320 96.900 135.120 97.200 ;
        RECT 137.820 96.900 139.620 97.200 ;
        RECT 133.320 96.600 134.520 96.900 ;
        RECT 138.420 96.600 139.620 96.900 ;
        RECT 133.320 96.300 134.220 96.600 ;
        RECT 138.720 96.300 139.620 96.600 ;
        RECT 133.620 96.000 133.920 96.300 ;
        RECT 135.420 96.000 135.720 96.300 ;
        RECT 136.020 96.000 136.320 96.300 ;
        RECT 136.620 96.000 136.920 96.300 ;
        RECT 137.220 96.000 137.520 96.300 ;
        RECT 139.020 96.000 139.320 96.300 ;
        RECT 135.420 95.400 137.520 96.000 ;
        RECT 134.820 95.100 136.020 95.400 ;
        RECT 136.920 95.100 137.820 95.400 ;
        RECT 134.820 94.800 136.320 95.100 ;
        RECT 136.620 94.800 138.420 95.100 ;
        RECT 134.520 94.500 135.120 94.800 ;
        RECT 135.720 94.500 137.220 94.800 ;
        RECT 137.820 94.500 138.420 94.800 ;
        RECT 134.520 94.200 134.820 94.500 ;
        RECT 134.220 93.900 134.820 94.200 ;
        RECT 134.220 93.600 135.120 93.900 ;
        RECT 136.020 93.600 136.920 94.500 ;
        RECT 138.120 94.200 138.420 94.500 ;
        RECT 138.120 93.900 138.720 94.200 ;
        RECT 137.820 93.600 138.720 93.900 ;
        RECT 134.220 92.400 138.720 93.600 ;
        RECT 134.520 91.800 138.420 92.400 ;
        RECT 135.120 91.500 137.820 91.800 ;
        RECT 138.610 91.760 140.000 92.200 ;
        RECT 139.440 91.590 140.000 91.760 ;
        RECT 135.120 91.200 137.520 91.500 ;
        RECT 23.740 89.150 24.940 89.450 ;
        RECT 25.240 89.150 26.440 89.450 ;
        RECT 28.060 89.350 29.120 89.560 ;
        RECT 21.940 88.850 24.340 89.150 ;
        RECT 25.840 88.850 27.940 89.150 ;
        RECT 21.940 88.550 23.740 88.850 ;
        RECT 26.440 88.550 28.240 88.850 ;
        RECT 21.940 88.250 23.140 88.550 ;
        RECT 27.040 88.250 28.240 88.550 ;
        RECT 21.940 87.950 22.840 88.250 ;
        RECT 27.340 87.950 28.240 88.250 ;
        RECT 22.240 87.650 22.540 87.950 ;
        RECT 24.040 87.650 24.340 87.950 ;
        RECT 24.640 87.650 24.940 87.950 ;
        RECT 25.240 87.650 25.540 87.950 ;
        RECT 25.840 87.650 26.140 87.950 ;
        RECT 27.640 87.650 27.940 87.950 ;
        RECT 24.040 87.050 26.140 87.650 ;
        RECT 23.440 86.750 24.640 87.050 ;
        RECT 25.540 86.750 26.440 87.050 ;
        RECT 23.440 86.450 24.940 86.750 ;
        RECT 25.240 86.450 27.040 86.750 ;
        RECT 23.140 86.150 23.740 86.450 ;
        RECT 24.340 86.150 25.840 86.450 ;
        RECT 26.440 86.150 27.040 86.450 ;
        RECT 23.140 85.850 23.440 86.150 ;
        RECT 22.840 85.550 23.440 85.850 ;
        RECT 22.840 85.250 23.740 85.550 ;
        RECT 24.640 85.250 25.540 86.150 ;
        RECT 26.740 85.850 27.040 86.150 ;
        RECT 26.740 85.550 27.340 85.850 ;
        RECT 26.440 85.250 27.340 85.550 ;
        RECT 22.840 84.050 27.340 85.250 ;
        RECT 23.140 83.450 27.040 84.050 ;
        RECT 23.740 83.150 26.440 83.450 ;
        RECT 27.230 83.410 28.620 83.850 ;
        RECT 28.060 83.240 28.620 83.410 ;
        RECT 23.740 82.850 26.140 83.150 ;
        RECT 30.520 73.030 31.020 89.560 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 131.830 89.560 133.240 90.060 ;
        RECT 127.360 88.590 129.760 88.890 ;
        RECT 127.360 88.290 130.060 88.590 ;
        RECT 131.790 88.320 132.240 88.430 ;
        RECT 126.760 87.690 130.660 88.290 ;
        RECT 131.130 87.820 132.240 88.320 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 126.460 86.490 130.960 87.690 ;
        RECT 126.460 86.190 127.360 86.490 ;
        RECT 126.460 85.890 127.060 86.190 ;
        RECT 126.760 85.590 127.060 85.890 ;
        RECT 128.260 85.590 129.160 86.490 ;
        RECT 130.060 86.190 130.960 86.490 ;
        RECT 130.360 85.890 130.960 86.190 ;
        RECT 130.360 85.590 130.660 85.890 ;
        RECT 126.760 85.290 127.360 85.590 ;
        RECT 127.960 85.290 129.460 85.590 ;
        RECT 130.060 85.290 130.660 85.590 ;
        RECT 127.060 84.990 128.560 85.290 ;
        RECT 128.860 84.990 130.660 85.290 ;
        RECT 127.060 84.690 128.260 84.990 ;
        RECT 129.160 84.690 130.060 84.990 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
        RECT 127.660 84.090 129.760 84.690 ;
        RECT 125.860 83.790 126.760 84.090 ;
        RECT 127.660 83.790 127.960 84.090 ;
        RECT 128.260 83.790 128.560 84.090 ;
        RECT 128.860 83.790 129.160 84.090 ;
        RECT 129.460 83.790 129.760 84.090 ;
        RECT 130.660 83.790 131.560 84.090 ;
        RECT 125.560 83.190 127.060 83.790 ;
        RECT 130.360 83.190 131.860 83.790 ;
        RECT 125.860 82.890 127.660 83.190 ;
        RECT 129.760 82.890 131.560 83.190 ;
        RECT 126.760 82.590 127.960 82.890 ;
        RECT 129.460 82.590 130.660 82.890 ;
        RECT 132.740 82.590 133.240 89.560 ;
        RECT 124.460 82.320 125.570 82.590 ;
        RECT 33.810 79.230 36.210 79.530 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 122.380 81.820 125.570 82.320 ;
        RECT 127.360 82.290 128.560 82.590 ;
        RECT 128.860 82.290 130.060 82.590 ;
        RECT 33.810 78.930 36.510 79.230 ;
        RECT 38.130 78.970 38.690 79.140 ;
        RECT 33.210 78.330 37.110 78.930 ;
        RECT 37.300 78.530 38.690 78.970 ;
        RECT 32.910 77.130 37.410 78.330 ;
        RECT 32.910 76.830 33.810 77.130 ;
        RECT 32.910 76.530 33.510 76.830 ;
        RECT 33.210 76.230 33.510 76.530 ;
        RECT 34.710 76.230 35.610 77.130 ;
        RECT 36.510 76.830 37.410 77.130 ;
        RECT 36.810 76.530 37.410 76.830 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
        RECT 36.810 76.230 37.110 76.530 ;
        RECT 33.210 75.930 33.810 76.230 ;
        RECT 34.410 75.930 35.910 76.230 ;
        RECT 36.510 75.930 37.110 76.230 ;
        RECT 33.510 75.630 35.010 75.930 ;
        RECT 35.310 75.630 37.110 75.930 ;
        RECT 33.510 75.330 34.710 75.630 ;
        RECT 35.610 75.330 36.510 75.630 ;
        RECT 34.110 74.730 36.210 75.330 ;
        RECT 32.310 74.430 32.610 74.730 ;
        RECT 34.110 74.430 34.410 74.730 ;
        RECT 34.710 74.430 35.010 74.730 ;
        RECT 35.310 74.430 35.610 74.730 ;
        RECT 35.910 74.430 36.210 74.730 ;
        RECT 37.710 74.430 38.010 74.730 ;
        RECT 32.010 74.130 32.910 74.430 ;
        RECT 37.410 74.130 38.310 74.430 ;
        RECT 32.010 73.830 33.210 74.130 ;
        RECT 37.110 73.830 38.310 74.130 ;
        RECT 32.010 73.530 33.810 73.830 ;
        RECT 36.510 73.530 38.310 73.830 ;
        RECT 32.010 73.230 34.410 73.530 ;
        RECT 35.910 73.230 38.010 73.530 ;
        RECT 30.520 72.300 32.020 73.030 ;
        RECT 33.810 72.930 35.010 73.230 ;
        RECT 35.310 72.930 36.510 73.230 ;
        RECT 115.190 73.140 117.590 73.440 ;
        RECT 34.410 72.330 35.910 72.930 ;
        RECT 38.130 72.800 39.190 73.030 ;
        RECT 115.190 72.840 117.890 73.140 ;
        RECT 119.510 72.880 120.070 73.050 ;
        RECT 30.910 72.030 32.020 72.300 ;
        RECT 33.810 72.030 35.010 72.330 ;
        RECT 35.310 72.030 36.510 72.330 ;
        RECT 38.130 72.300 41.210 72.800 ;
        RECT 38.130 72.030 39.190 72.300 ;
        RECT 33.210 71.730 34.410 72.030 ;
        RECT 35.910 71.730 37.110 72.030 ;
        RECT 32.310 71.430 34.110 71.730 ;
        RECT 36.210 71.430 38.010 71.730 ;
        RECT 32.010 70.830 33.510 71.430 ;
        RECT 36.810 70.830 38.310 71.430 ;
        RECT 32.310 70.530 33.210 70.830 ;
        RECT 34.110 70.530 34.410 70.830 ;
        RECT 34.710 70.530 35.010 70.830 ;
        RECT 35.310 70.530 35.610 70.830 ;
        RECT 35.910 70.530 36.210 70.830 ;
        RECT 37.110 70.530 38.010 70.830 ;
        RECT 34.110 69.930 36.210 70.530 ;
        RECT 33.510 69.630 34.710 69.930 ;
        RECT 35.610 69.630 36.510 69.930 ;
        RECT 33.510 69.330 35.010 69.630 ;
        RECT 35.310 69.330 37.110 69.630 ;
        RECT 33.210 69.030 33.810 69.330 ;
        RECT 34.410 69.030 35.910 69.330 ;
        RECT 36.510 69.030 37.110 69.330 ;
        RECT 33.210 68.730 33.510 69.030 ;
        RECT 32.910 68.430 33.510 68.730 ;
        RECT 32.910 68.130 33.810 68.430 ;
        RECT 34.710 68.130 35.610 69.030 ;
        RECT 36.810 68.730 37.110 69.030 ;
        RECT 36.810 68.430 37.410 68.730 ;
        RECT 36.510 68.130 37.410 68.430 ;
        RECT 32.910 66.930 37.410 68.130 ;
        RECT 33.210 66.330 37.110 66.930 ;
        RECT 33.810 66.030 36.510 66.330 ;
        RECT 37.580 66.300 38.690 66.800 ;
        RECT 38.240 66.190 38.690 66.300 ;
        RECT 33.810 65.730 36.210 66.030 ;
        RECT 40.710 61.630 41.210 72.300 ;
        RECT 114.590 72.240 118.490 72.840 ;
        RECT 118.680 72.440 120.070 72.880 ;
        RECT 114.290 71.040 118.790 72.240 ;
        RECT 114.290 70.740 115.190 71.040 ;
        RECT 114.290 70.440 114.890 70.740 ;
        RECT 114.590 70.140 114.890 70.440 ;
        RECT 116.090 70.140 116.990 71.040 ;
        RECT 117.890 70.740 118.790 71.040 ;
        RECT 118.190 70.440 118.790 70.740 ;
        RECT 118.190 70.140 118.490 70.440 ;
        RECT 114.590 69.840 115.190 70.140 ;
        RECT 115.790 69.840 117.290 70.140 ;
        RECT 117.890 69.840 118.490 70.140 ;
        RECT 114.890 69.540 116.390 69.840 ;
        RECT 116.690 69.540 118.490 69.840 ;
        RECT 114.890 69.240 116.090 69.540 ;
        RECT 116.990 69.240 117.890 69.540 ;
        RECT 115.490 68.640 117.590 69.240 ;
        RECT 47.790 68.080 50.190 68.380 ;
        RECT 113.690 68.340 113.990 68.640 ;
        RECT 115.490 68.340 115.790 68.640 ;
        RECT 116.090 68.340 116.390 68.640 ;
        RECT 116.690 68.340 116.990 68.640 ;
        RECT 117.290 68.340 117.590 68.640 ;
        RECT 119.090 68.340 119.390 68.640 ;
        RECT 47.790 67.780 50.490 68.080 ;
        RECT 113.390 68.040 114.290 68.340 ;
        RECT 118.790 68.040 119.690 68.340 ;
        RECT 52.110 67.820 52.670 67.990 ;
        RECT 47.190 67.180 51.090 67.780 ;
        RECT 51.280 67.380 52.670 67.820 ;
        RECT 113.390 67.740 114.590 68.040 ;
        RECT 118.490 67.740 119.690 68.040 ;
        RECT 113.390 67.440 115.190 67.740 ;
        RECT 117.890 67.440 119.690 67.740 ;
        RECT 46.890 65.980 51.390 67.180 ;
        RECT 113.390 67.140 115.790 67.440 ;
        RECT 117.290 67.140 119.390 67.440 ;
        RECT 112.290 66.710 113.400 66.940 ;
        RECT 115.190 66.840 116.390 67.140 ;
        RECT 116.690 66.840 117.890 67.140 ;
        RECT 46.890 65.680 47.790 65.980 ;
        RECT 46.890 65.380 47.490 65.680 ;
        RECT 47.190 65.080 47.490 65.380 ;
        RECT 48.690 65.080 49.590 65.980 ;
        RECT 50.490 65.680 51.390 65.980 ;
        RECT 50.790 65.380 51.390 65.680 ;
        RECT 111.900 65.940 113.400 66.710 ;
        RECT 115.790 66.240 117.290 66.840 ;
        RECT 119.510 66.710 120.570 66.940 ;
        RECT 122.380 66.710 122.880 81.820 ;
        RECT 124.460 81.590 125.570 81.820 ;
        RECT 127.960 81.690 129.460 82.290 ;
        RECT 131.680 81.820 133.240 82.590 ;
        RECT 127.360 81.390 128.560 81.690 ;
        RECT 128.860 81.390 130.060 81.690 ;
        RECT 131.680 81.590 132.740 81.820 ;
        RECT 125.560 81.090 127.960 81.390 ;
        RECT 129.460 81.090 131.560 81.390 ;
        RECT 125.560 80.790 127.360 81.090 ;
        RECT 130.060 80.790 131.860 81.090 ;
        RECT 125.560 80.490 126.760 80.790 ;
        RECT 130.660 80.490 131.860 80.790 ;
        RECT 125.560 80.190 126.460 80.490 ;
        RECT 130.960 80.190 131.860 80.490 ;
        RECT 125.860 79.890 126.160 80.190 ;
        RECT 127.660 79.890 127.960 80.190 ;
        RECT 128.260 79.890 128.560 80.190 ;
        RECT 128.860 79.890 129.160 80.190 ;
        RECT 129.460 79.890 129.760 80.190 ;
        RECT 131.260 79.890 131.560 80.190 ;
        RECT 127.660 79.290 129.760 79.890 ;
        RECT 127.060 78.990 128.260 79.290 ;
        RECT 129.160 78.990 130.060 79.290 ;
        RECT 127.060 78.690 128.560 78.990 ;
        RECT 128.860 78.690 130.660 78.990 ;
        RECT 126.760 78.390 127.360 78.690 ;
        RECT 127.960 78.390 129.460 78.690 ;
        RECT 130.060 78.390 130.660 78.690 ;
        RECT 126.760 78.090 127.060 78.390 ;
        RECT 126.460 77.790 127.060 78.090 ;
        RECT 126.460 77.490 127.360 77.790 ;
        RECT 128.260 77.490 129.160 78.390 ;
        RECT 130.360 78.090 130.660 78.390 ;
        RECT 130.360 77.790 130.960 78.090 ;
        RECT 130.060 77.490 130.960 77.790 ;
        RECT 126.460 76.290 130.960 77.490 ;
        RECT 126.760 75.690 130.660 76.290 ;
        RECT 127.360 75.390 130.060 75.690 ;
        RECT 130.850 75.650 132.240 76.090 ;
        RECT 131.680 75.480 132.240 75.650 ;
        RECT 127.360 75.090 129.760 75.390 ;
        RECT 115.190 65.940 116.390 66.240 ;
        RECT 116.690 65.940 117.890 66.240 ;
        RECT 119.510 66.210 122.880 66.710 ;
        RECT 119.510 65.940 120.570 66.210 ;
        RECT 50.790 65.080 51.090 65.380 ;
        RECT 47.190 64.780 47.790 65.080 ;
        RECT 48.390 64.780 49.890 65.080 ;
        RECT 50.490 64.780 51.090 65.080 ;
        RECT 47.490 64.480 48.990 64.780 ;
        RECT 49.290 64.480 51.090 64.780 ;
        RECT 47.490 64.180 48.690 64.480 ;
        RECT 49.590 64.180 50.490 64.480 ;
        RECT 99.710 64.190 102.110 64.490 ;
        RECT 48.090 63.580 50.190 64.180 ;
        RECT 99.710 63.890 102.410 64.190 ;
        RECT 104.030 63.930 104.590 64.100 ;
        RECT 46.290 63.280 46.590 63.580 ;
        RECT 48.090 63.280 48.390 63.580 ;
        RECT 48.690 63.280 48.990 63.580 ;
        RECT 49.290 63.280 49.590 63.580 ;
        RECT 49.890 63.280 50.190 63.580 ;
        RECT 51.690 63.280 51.990 63.580 ;
        RECT 99.110 63.290 103.010 63.890 ;
        RECT 103.200 63.490 104.590 63.930 ;
        RECT 45.990 62.980 46.890 63.280 ;
        RECT 51.390 62.980 52.290 63.280 ;
        RECT 45.990 62.680 47.190 62.980 ;
        RECT 51.090 62.680 52.290 62.980 ;
        RECT 45.990 62.380 47.790 62.680 ;
        RECT 50.490 62.380 52.290 62.680 ;
        RECT 45.990 62.080 48.390 62.380 ;
        RECT 49.890 62.080 51.990 62.380 ;
        RECT 98.810 62.090 103.310 63.290 ;
        RECT 44.890 61.650 46.000 61.880 ;
        RECT 47.790 61.780 48.990 62.080 ;
        RECT 49.290 61.780 50.490 62.080 ;
        RECT 44.500 61.630 46.000 61.650 ;
        RECT 40.710 61.130 46.000 61.630 ;
        RECT 48.390 61.180 49.890 61.780 ;
        RECT 52.110 61.650 53.170 61.880 ;
        RECT 44.890 60.880 46.000 61.130 ;
        RECT 47.790 60.880 48.990 61.180 ;
        RECT 49.290 60.880 50.490 61.180 ;
        RECT 52.110 61.150 57.830 61.650 ;
        RECT 64.440 61.550 66.840 61.850 ;
        RECT 98.810 61.790 99.710 62.090 ;
        RECT 64.440 61.250 67.140 61.550 ;
        RECT 98.810 61.490 99.410 61.790 ;
        RECT 68.760 61.290 69.320 61.460 ;
        RECT 52.110 60.880 53.170 61.150 ;
        RECT 47.190 60.580 48.390 60.880 ;
        RECT 49.890 60.580 51.090 60.880 ;
        RECT 46.290 60.280 48.090 60.580 ;
        RECT 50.190 60.280 51.990 60.580 ;
        RECT 45.990 59.680 47.490 60.280 ;
        RECT 50.790 59.680 52.290 60.280 ;
        RECT 46.290 59.380 47.190 59.680 ;
        RECT 48.090 59.380 48.390 59.680 ;
        RECT 48.690 59.380 48.990 59.680 ;
        RECT 49.290 59.380 49.590 59.680 ;
        RECT 49.890 59.380 50.190 59.680 ;
        RECT 51.090 59.380 51.990 59.680 ;
        RECT 48.090 58.780 50.190 59.380 ;
        RECT 47.490 58.480 48.690 58.780 ;
        RECT 49.590 58.480 50.490 58.780 ;
        RECT 47.490 58.180 48.990 58.480 ;
        RECT 49.290 58.180 51.090 58.480 ;
        RECT 47.190 57.880 47.790 58.180 ;
        RECT 48.390 57.880 49.890 58.180 ;
        RECT 50.490 57.880 51.090 58.180 ;
        RECT 47.190 57.580 47.490 57.880 ;
        RECT 46.890 57.280 47.490 57.580 ;
        RECT 46.890 56.980 47.790 57.280 ;
        RECT 48.690 56.980 49.590 57.880 ;
        RECT 50.790 57.580 51.090 57.880 ;
        RECT 50.790 57.280 51.390 57.580 ;
        RECT 50.490 56.980 51.390 57.280 ;
        RECT 46.890 55.780 51.390 56.980 ;
        RECT 47.190 55.180 51.090 55.780 ;
        RECT 47.790 54.880 50.490 55.180 ;
        RECT 51.560 55.150 52.670 55.650 ;
        RECT 52.220 55.040 52.670 55.150 ;
        RECT 57.330 55.140 57.830 61.150 ;
        RECT 63.840 60.650 67.740 61.250 ;
        RECT 67.930 60.850 69.320 61.290 ;
        RECT 99.110 61.190 99.410 61.490 ;
        RECT 100.610 61.190 101.510 62.090 ;
        RECT 102.410 61.790 103.310 62.090 ;
        RECT 102.710 61.490 103.310 61.790 ;
        RECT 102.710 61.190 103.010 61.490 ;
        RECT 99.110 60.890 99.710 61.190 ;
        RECT 100.310 60.890 101.810 61.190 ;
        RECT 102.410 60.890 103.010 61.190 ;
        RECT 63.540 59.450 68.040 60.650 ;
        RECT 99.410 60.590 100.910 60.890 ;
        RECT 101.210 60.590 103.010 60.890 ;
        RECT 82.270 60.210 84.670 60.510 ;
        RECT 99.410 60.290 100.610 60.590 ;
        RECT 101.510 60.290 102.410 60.590 ;
        RECT 82.270 59.910 84.970 60.210 ;
        RECT 86.590 59.950 87.150 60.120 ;
        RECT 63.540 59.150 64.440 59.450 ;
        RECT 63.540 58.850 64.140 59.150 ;
        RECT 63.840 58.550 64.140 58.850 ;
        RECT 65.340 58.550 66.240 59.450 ;
        RECT 67.140 59.150 68.040 59.450 ;
        RECT 81.670 59.310 85.570 59.910 ;
        RECT 85.760 59.510 87.150 59.950 ;
        RECT 100.010 59.690 102.110 60.290 ;
        RECT 98.210 59.390 98.510 59.690 ;
        RECT 100.010 59.390 100.310 59.690 ;
        RECT 100.610 59.390 100.910 59.690 ;
        RECT 101.210 59.390 101.510 59.690 ;
        RECT 101.810 59.390 102.110 59.690 ;
        RECT 103.610 59.390 103.910 59.690 ;
        RECT 67.440 58.850 68.040 59.150 ;
        RECT 67.440 58.550 67.740 58.850 ;
        RECT 63.840 58.250 64.440 58.550 ;
        RECT 65.040 58.250 66.540 58.550 ;
        RECT 67.140 58.250 67.740 58.550 ;
        RECT 64.140 57.950 65.640 58.250 ;
        RECT 65.940 57.950 67.740 58.250 ;
        RECT 81.370 58.110 85.870 59.310 ;
        RECT 97.910 59.090 98.810 59.390 ;
        RECT 103.310 59.090 104.210 59.390 ;
        RECT 97.910 58.790 99.110 59.090 ;
        RECT 103.010 58.790 104.210 59.090 ;
        RECT 97.910 58.490 99.710 58.790 ;
        RECT 102.410 58.490 104.210 58.790 ;
        RECT 97.910 58.190 100.310 58.490 ;
        RECT 101.810 58.190 103.910 58.490 ;
        RECT 64.140 57.650 65.340 57.950 ;
        RECT 66.240 57.650 67.140 57.950 ;
        RECT 81.370 57.810 82.270 58.110 ;
        RECT 64.740 57.050 66.840 57.650 ;
        RECT 81.370 57.510 81.970 57.810 ;
        RECT 81.670 57.210 81.970 57.510 ;
        RECT 83.170 57.210 84.070 58.110 ;
        RECT 84.970 57.810 85.870 58.110 ;
        RECT 85.270 57.510 85.870 57.810 ;
        RECT 96.810 57.760 97.920 57.990 ;
        RECT 99.710 57.890 100.910 58.190 ;
        RECT 101.210 57.890 102.410 58.190 ;
        RECT 85.270 57.210 85.570 57.510 ;
        RECT 96.420 57.260 97.920 57.760 ;
        RECT 100.310 57.290 101.810 57.890 ;
        RECT 104.030 57.760 105.090 57.990 ;
        RECT 104.030 57.730 105.590 57.760 ;
        RECT 111.900 57.730 112.400 65.940 ;
        RECT 114.590 65.640 115.790 65.940 ;
        RECT 117.290 65.640 118.490 65.940 ;
        RECT 113.690 65.340 115.490 65.640 ;
        RECT 117.590 65.340 119.390 65.640 ;
        RECT 113.390 64.740 114.890 65.340 ;
        RECT 118.190 64.740 119.690 65.340 ;
        RECT 113.690 64.440 114.590 64.740 ;
        RECT 115.490 64.440 115.790 64.740 ;
        RECT 116.090 64.440 116.390 64.740 ;
        RECT 116.690 64.440 116.990 64.740 ;
        RECT 117.290 64.440 117.590 64.740 ;
        RECT 118.490 64.440 119.390 64.740 ;
        RECT 115.490 63.840 117.590 64.440 ;
        RECT 114.890 63.540 116.090 63.840 ;
        RECT 116.990 63.540 117.890 63.840 ;
        RECT 114.890 63.240 116.390 63.540 ;
        RECT 116.690 63.240 118.490 63.540 ;
        RECT 114.590 62.940 115.190 63.240 ;
        RECT 115.790 62.940 117.290 63.240 ;
        RECT 117.890 62.940 118.490 63.240 ;
        RECT 114.590 62.640 114.890 62.940 ;
        RECT 114.290 62.340 114.890 62.640 ;
        RECT 114.290 62.040 115.190 62.340 ;
        RECT 116.090 62.040 116.990 62.940 ;
        RECT 118.190 62.640 118.490 62.940 ;
        RECT 118.190 62.340 118.790 62.640 ;
        RECT 117.890 62.040 118.790 62.340 ;
        RECT 114.290 60.840 118.790 62.040 ;
        RECT 114.590 60.240 118.490 60.840 ;
        RECT 115.190 59.940 117.890 60.240 ;
        RECT 118.960 60.210 120.070 60.710 ;
        RECT 119.620 60.100 120.070 60.210 ;
        RECT 115.190 59.640 117.590 59.940 ;
        RECT 62.940 56.750 63.240 57.050 ;
        RECT 64.740 56.750 65.040 57.050 ;
        RECT 65.340 56.750 65.640 57.050 ;
        RECT 65.940 56.750 66.240 57.050 ;
        RECT 66.540 56.750 66.840 57.050 ;
        RECT 68.340 56.750 68.640 57.050 ;
        RECT 81.670 56.910 82.270 57.210 ;
        RECT 82.870 56.910 84.370 57.210 ;
        RECT 84.970 56.910 85.570 57.210 ;
        RECT 62.640 56.450 63.540 56.750 ;
        RECT 68.040 56.450 68.940 56.750 ;
        RECT 62.640 56.150 63.840 56.450 ;
        RECT 67.740 56.150 68.940 56.450 ;
        RECT 81.970 56.610 83.470 56.910 ;
        RECT 83.770 56.610 85.570 56.910 ;
        RECT 96.430 56.990 97.920 57.260 ;
        RECT 99.710 56.990 100.910 57.290 ;
        RECT 101.210 56.990 102.410 57.290 ;
        RECT 104.030 57.230 112.400 57.730 ;
        RECT 104.030 56.990 105.090 57.230 ;
        RECT 81.970 56.310 83.170 56.610 ;
        RECT 84.070 56.310 84.970 56.610 ;
        RECT 62.640 55.850 64.440 56.150 ;
        RECT 67.140 55.850 68.940 56.150 ;
        RECT 62.640 55.550 65.040 55.850 ;
        RECT 66.540 55.550 68.640 55.850 ;
        RECT 82.570 55.710 84.670 56.310 ;
        RECT 61.540 55.140 62.650 55.350 ;
        RECT 64.440 55.250 65.640 55.550 ;
        RECT 65.940 55.250 67.140 55.550 ;
        RECT 80.770 55.410 81.070 55.710 ;
        RECT 82.570 55.410 82.870 55.710 ;
        RECT 83.170 55.410 83.470 55.710 ;
        RECT 83.770 55.410 84.070 55.710 ;
        RECT 84.370 55.410 84.670 55.710 ;
        RECT 86.170 55.410 86.470 55.710 ;
        RECT 47.790 54.580 50.190 54.880 ;
        RECT 57.330 54.640 62.650 55.140 ;
        RECT 65.040 54.650 66.540 55.250 ;
        RECT 68.760 55.120 69.820 55.350 ;
        RECT 61.150 54.620 62.650 54.640 ;
        RECT 61.540 54.350 62.650 54.620 ;
        RECT 64.440 54.350 65.640 54.650 ;
        RECT 65.940 54.350 67.140 54.650 ;
        RECT 68.760 54.620 74.620 55.120 ;
        RECT 68.760 54.350 69.820 54.620 ;
        RECT 63.840 54.050 65.040 54.350 ;
        RECT 66.540 54.050 67.740 54.350 ;
        RECT 62.940 53.750 64.740 54.050 ;
        RECT 66.840 53.750 68.640 54.050 ;
        RECT 74.120 53.750 74.620 54.620 ;
        RECT 80.470 55.110 81.370 55.410 ;
        RECT 85.870 55.110 86.770 55.410 ;
        RECT 80.470 54.810 81.670 55.110 ;
        RECT 85.570 54.810 86.770 55.110 ;
        RECT 80.470 54.510 82.270 54.810 ;
        RECT 84.970 54.510 86.770 54.810 ;
        RECT 80.470 54.210 82.870 54.510 ;
        RECT 84.370 54.210 86.470 54.510 ;
        RECT 79.370 53.780 80.480 54.010 ;
        RECT 82.270 53.910 83.470 54.210 ;
        RECT 83.770 53.910 84.970 54.210 ;
        RECT 78.980 53.750 80.480 53.780 ;
        RECT 62.640 53.150 64.140 53.750 ;
        RECT 67.440 53.150 68.940 53.750 ;
        RECT 74.120 53.250 80.480 53.750 ;
        RECT 82.870 53.310 84.370 53.910 ;
        RECT 86.590 53.780 87.650 54.010 ;
        RECT 96.430 53.780 96.930 56.990 ;
        RECT 99.110 56.690 100.310 56.990 ;
        RECT 101.810 56.690 103.010 56.990 ;
        RECT 98.210 56.390 100.010 56.690 ;
        RECT 102.110 56.390 103.910 56.690 ;
        RECT 97.910 55.790 99.410 56.390 ;
        RECT 102.710 55.790 104.210 56.390 ;
        RECT 98.210 55.490 99.110 55.790 ;
        RECT 100.010 55.490 100.310 55.790 ;
        RECT 100.610 55.490 100.910 55.790 ;
        RECT 101.210 55.490 101.510 55.790 ;
        RECT 101.810 55.490 102.110 55.790 ;
        RECT 103.010 55.490 103.910 55.790 ;
        RECT 100.010 54.890 102.110 55.490 ;
        RECT 99.410 54.590 100.610 54.890 ;
        RECT 101.510 54.590 102.410 54.890 ;
        RECT 99.410 54.290 100.910 54.590 ;
        RECT 101.210 54.290 103.010 54.590 ;
        RECT 62.940 52.850 63.840 53.150 ;
        RECT 64.740 52.850 65.040 53.150 ;
        RECT 65.340 52.850 65.640 53.150 ;
        RECT 65.940 52.850 66.240 53.150 ;
        RECT 66.540 52.850 66.840 53.150 ;
        RECT 67.740 52.850 68.640 53.150 ;
        RECT 79.370 53.010 80.480 53.250 ;
        RECT 82.270 53.010 83.470 53.310 ;
        RECT 83.770 53.010 84.970 53.310 ;
        RECT 86.590 53.280 96.930 53.780 ;
        RECT 99.110 53.990 99.710 54.290 ;
        RECT 100.310 53.990 101.810 54.290 ;
        RECT 102.410 53.990 103.010 54.290 ;
        RECT 99.110 53.690 99.410 53.990 ;
        RECT 98.810 53.390 99.410 53.690 ;
        RECT 86.590 53.010 87.650 53.280 ;
        RECT 98.810 53.090 99.710 53.390 ;
        RECT 100.610 53.090 101.510 53.990 ;
        RECT 102.710 53.690 103.010 53.990 ;
        RECT 102.710 53.390 103.310 53.690 ;
        RECT 102.410 53.090 103.310 53.390 ;
        RECT 64.740 52.250 66.840 52.850 ;
        RECT 81.670 52.710 82.870 53.010 ;
        RECT 84.370 52.710 85.570 53.010 ;
        RECT 80.770 52.410 82.570 52.710 ;
        RECT 84.670 52.410 86.470 52.710 ;
        RECT 64.140 51.950 65.340 52.250 ;
        RECT 66.240 51.950 67.140 52.250 ;
        RECT 64.140 51.650 65.640 51.950 ;
        RECT 65.940 51.650 67.740 51.950 ;
        RECT 80.470 51.810 81.970 52.410 ;
        RECT 85.270 51.810 86.770 52.410 ;
        RECT 98.810 51.890 103.310 53.090 ;
        RECT 63.840 51.350 64.440 51.650 ;
        RECT 65.040 51.350 66.540 51.650 ;
        RECT 67.140 51.350 67.740 51.650 ;
        RECT 80.770 51.510 81.670 51.810 ;
        RECT 82.570 51.510 82.870 51.810 ;
        RECT 83.170 51.510 83.470 51.810 ;
        RECT 83.770 51.510 84.070 51.810 ;
        RECT 84.370 51.510 84.670 51.810 ;
        RECT 85.570 51.510 86.470 51.810 ;
        RECT 63.840 51.050 64.140 51.350 ;
        RECT 63.540 50.750 64.140 51.050 ;
        RECT 63.540 50.450 64.440 50.750 ;
        RECT 65.340 50.450 66.240 51.350 ;
        RECT 67.440 51.050 67.740 51.350 ;
        RECT 67.440 50.750 68.040 51.050 ;
        RECT 82.570 50.910 84.670 51.510 ;
        RECT 99.110 51.290 103.010 51.890 ;
        RECT 99.710 50.990 102.410 51.290 ;
        RECT 103.480 51.260 104.590 51.760 ;
        RECT 104.140 51.150 104.590 51.260 ;
        RECT 67.140 50.450 68.040 50.750 ;
        RECT 63.540 49.250 68.040 50.450 ;
        RECT 81.970 50.610 83.170 50.910 ;
        RECT 84.070 50.610 84.970 50.910 ;
        RECT 99.710 50.690 102.110 50.990 ;
        RECT 81.970 50.310 83.470 50.610 ;
        RECT 83.770 50.310 85.570 50.610 ;
        RECT 81.670 50.010 82.270 50.310 ;
        RECT 82.870 50.010 84.370 50.310 ;
        RECT 84.970 50.010 85.570 50.310 ;
        RECT 81.670 49.710 81.970 50.010 ;
        RECT 81.370 49.410 81.970 49.710 ;
        RECT 63.840 48.650 67.740 49.250 ;
        RECT 64.440 48.350 67.140 48.650 ;
        RECT 68.210 48.620 69.320 49.120 ;
        RECT 68.870 48.510 69.320 48.620 ;
        RECT 81.370 49.110 82.270 49.410 ;
        RECT 83.170 49.110 84.070 50.010 ;
        RECT 85.270 49.710 85.570 50.010 ;
        RECT 85.270 49.410 85.870 49.710 ;
        RECT 84.970 49.110 85.870 49.410 ;
        RECT 64.440 48.050 66.840 48.350 ;
        RECT 81.370 47.910 85.870 49.110 ;
        RECT 81.670 47.310 85.570 47.910 ;
        RECT 82.270 47.010 84.970 47.310 ;
        RECT 86.040 47.280 87.150 47.780 ;
        RECT 86.700 47.170 87.150 47.280 ;
        RECT 82.270 46.710 84.670 47.010 ;
      LAYER met2 ;
        RECT 85.860 223.640 86.180 224.140 ;
        RECT 88.620 223.640 88.940 224.140 ;
        RECT 85.870 222.770 86.130 223.640 ;
        RECT 64.330 222.510 86.130 222.770 ;
        RECT 64.330 219.110 64.590 222.510 ;
        RECT 88.640 222.250 88.900 223.640 ;
        RECT 74.040 221.990 88.900 222.250 ;
        RECT 64.320 218.750 64.630 219.110 ;
        RECT 74.040 219.070 74.300 221.990 ;
        RECT 91.380 221.830 91.700 224.140 ;
        RECT 83.680 221.570 91.700 221.830 ;
        RECT 83.680 219.170 83.940 221.570 ;
        RECT 91.770 220.815 92.250 221.395 ;
        RECT 90.300 219.355 90.760 220.010 ;
        RECT 61.410 218.030 62.100 218.730 ;
        RECT 73.990 218.710 74.300 219.070 ;
        RECT 83.630 218.810 83.940 219.170 ;
        RECT 60.100 215.395 60.650 215.775 ;
        RECT 52.200 215.130 52.700 215.235 ;
        RECT 67.210 215.130 67.770 216.740 ;
        RECT 52.200 214.680 54.650 215.130 ;
        RECT 52.200 214.635 52.700 214.680 ;
        RECT 58.680 214.450 59.280 214.750 ;
        RECT 61.380 214.450 62.280 214.750 ;
        RECT 66.380 214.570 67.770 215.130 ;
        RECT 54.780 213.550 56.580 213.850 ;
        RECT 58.380 213.550 59.580 214.450 ;
        RECT 61.080 214.150 62.580 214.450 ;
        RECT 61.080 213.850 62.280 214.150 ;
        RECT 61.080 213.550 61.980 213.850 ;
        RECT 64.380 213.550 66.180 213.850 ;
        RECT 54.180 213.250 57.480 213.550 ;
        RECT 58.680 213.250 59.880 213.550 ;
        RECT 54.180 212.950 56.280 213.250 ;
        RECT 56.880 212.950 57.480 213.250 ;
        RECT 59.280 212.950 59.880 213.250 ;
        RECT 61.080 212.950 61.680 213.550 ;
        RECT 63.480 213.250 66.780 213.550 ;
        RECT 63.480 212.950 64.080 213.250 ;
        RECT 64.680 212.950 66.780 213.250 ;
        RECT 53.880 212.650 55.980 212.950 ;
        RECT 53.580 212.050 55.980 212.650 ;
        RECT 57.180 212.650 57.780 212.950 ;
        RECT 59.280 212.650 60.180 212.950 ;
        RECT 57.180 212.350 58.680 212.650 ;
        RECT 59.580 212.350 60.180 212.650 ;
        RECT 60.780 212.350 61.380 212.950 ;
        RECT 63.180 212.650 63.780 212.950 ;
        RECT 62.280 212.350 63.780 212.650 ;
        RECT 64.980 212.650 67.080 212.950 ;
        RECT 56.880 212.050 58.380 212.350 ;
        RECT 53.580 211.750 57.480 212.050 ;
        RECT 57.780 211.750 58.680 212.050 ;
        RECT 59.880 211.750 61.080 212.350 ;
        RECT 62.580 212.050 64.080 212.350 ;
        RECT 64.980 212.050 67.380 212.650 ;
        RECT 62.280 211.750 63.180 212.050 ;
        RECT 63.480 211.750 67.380 212.050 ;
        RECT 53.580 211.450 57.180 211.750 ;
        RECT 57.780 211.450 58.380 211.750 ;
        RECT 60.180 211.450 60.780 211.750 ;
        RECT 62.580 211.450 63.180 211.750 ;
        RECT 63.780 211.450 67.380 211.750 ;
        RECT 53.580 211.150 57.480 211.450 ;
        RECT 57.780 211.150 58.680 211.450 ;
        RECT 53.580 210.250 55.980 211.150 ;
        RECT 56.880 210.850 58.380 211.150 ;
        RECT 59.880 210.850 61.080 211.450 ;
        RECT 62.280 211.150 63.180 211.450 ;
        RECT 63.480 211.150 67.380 211.450 ;
        RECT 62.580 210.850 64.080 211.150 ;
        RECT 57.180 210.550 58.680 210.850 ;
        RECT 59.580 210.550 60.180 210.850 ;
        RECT 57.180 210.250 57.780 210.550 ;
        RECT 54.180 209.950 56.280 210.250 ;
        RECT 56.880 209.950 57.780 210.250 ;
        RECT 59.280 210.250 60.180 210.550 ;
        RECT 60.780 210.250 61.380 210.850 ;
        RECT 62.280 210.550 63.780 210.850 ;
        RECT 63.180 210.250 63.780 210.550 ;
        RECT 64.980 210.250 67.380 211.150 ;
        RECT 59.280 209.950 59.880 210.250 ;
        RECT 54.180 209.650 57.180 209.950 ;
        RECT 58.680 209.650 59.880 209.950 ;
        RECT 61.080 209.650 61.680 210.250 ;
        RECT 63.180 209.950 64.080 210.250 ;
        RECT 64.680 209.950 66.780 210.250 ;
        RECT 63.780 209.650 66.780 209.950 ;
        RECT 54.780 209.350 56.580 209.650 ;
        RECT 58.380 208.750 59.580 209.650 ;
        RECT 61.080 209.350 61.980 209.650 ;
        RECT 64.380 209.350 66.180 209.650 ;
        RECT 61.080 209.050 62.280 209.350 ;
        RECT 61.080 208.750 62.580 209.050 ;
        RECT 58.680 208.450 59.280 208.750 ;
        RECT 61.080 208.450 62.280 208.750 ;
        RECT 79.445 187.600 81.440 187.610 ;
        RECT 78.540 187.585 82.340 187.600 ;
        RECT 77.635 187.555 83.245 187.585 ;
        RECT 76.730 187.515 84.150 187.555 ;
        RECT 75.825 187.465 85.055 187.515 ;
        RECT 74.920 187.405 85.960 187.465 ;
        RECT 74.020 187.330 86.860 187.405 ;
        RECT 73.115 187.245 87.765 187.330 ;
        RECT 72.215 187.150 88.665 187.245 ;
        RECT 71.315 187.040 89.565 187.150 ;
        RECT 70.420 186.920 90.460 187.040 ;
        RECT 69.520 186.790 91.360 186.920 ;
        RECT 68.625 186.650 92.255 186.790 ;
        RECT 67.735 186.495 93.145 186.650 ;
        RECT 66.840 186.330 94.040 186.495 ;
        RECT 65.950 186.155 94.930 186.330 ;
        RECT 65.065 185.970 95.815 186.155 ;
        RECT 64.180 185.775 96.700 185.970 ;
        RECT 63.295 185.600 97.585 185.775 ;
        RECT 63.295 185.585 79.635 185.600 ;
        RECT 81.245 185.585 97.585 185.600 ;
        RECT 63.295 185.565 78.730 185.585 ;
        RECT 62.415 185.555 78.730 185.565 ;
        RECT 82.150 185.565 97.585 185.585 ;
        RECT 82.150 185.555 98.465 185.565 ;
        RECT 62.415 185.515 77.825 185.555 ;
        RECT 82.690 185.515 98.465 185.555 ;
        RECT 62.415 185.465 76.920 185.515 ;
        RECT 62.415 185.405 76.020 185.465 ;
        RECT 62.415 185.345 75.115 185.405 ;
        RECT 61.535 185.330 75.115 185.345 ;
        RECT 61.535 185.245 74.215 185.330 ;
        RECT 61.535 185.150 73.315 185.245 ;
        RECT 61.535 185.115 72.420 185.150 ;
        RECT 60.660 185.040 72.420 185.115 ;
        RECT 60.660 184.920 71.520 185.040 ;
        RECT 60.660 184.875 70.625 184.920 ;
        RECT 59.790 184.790 70.625 184.875 ;
        RECT 59.790 184.650 69.735 184.790 ;
        RECT 59.790 184.620 68.840 184.650 ;
        RECT 58.920 184.495 68.840 184.620 ;
        RECT 58.920 184.360 67.950 184.495 ;
        RECT 58.055 184.330 67.950 184.360 ;
        RECT 58.055 184.155 67.065 184.330 ;
        RECT 58.055 184.085 66.180 184.155 ;
        RECT 57.195 183.970 66.180 184.085 ;
        RECT 57.195 183.800 65.310 183.970 ;
        RECT 56.335 183.775 65.310 183.800 ;
        RECT 56.335 183.565 64.415 183.775 ;
        RECT 56.335 183.505 63.535 183.565 ;
        RECT 55.480 183.345 63.535 183.505 ;
        RECT 55.480 183.195 62.660 183.345 ;
        RECT 54.630 183.115 62.660 183.195 ;
        RECT 54.630 182.880 61.790 183.115 ;
        RECT 53.780 182.875 61.790 182.880 ;
        RECT 53.780 182.620 60.920 182.875 ;
        RECT 53.780 182.550 60.055 182.620 ;
        RECT 52.940 182.360 60.055 182.550 ;
        RECT 52.940 182.215 59.195 182.360 ;
        RECT 52.100 182.085 59.195 182.215 ;
        RECT 52.100 181.865 58.335 182.085 ;
        RECT 51.265 181.800 58.335 181.865 ;
        RECT 51.265 181.505 57.480 181.800 ;
        RECT 50.435 181.195 56.630 181.505 ;
        RECT 50.435 181.135 55.780 181.195 ;
        RECT 49.605 180.880 55.780 181.135 ;
        RECT 49.605 180.755 54.940 180.880 ;
        RECT 48.785 180.550 54.940 180.755 ;
        RECT 48.785 180.365 54.100 180.550 ;
        RECT 47.970 180.215 54.100 180.365 ;
        RECT 47.970 179.965 53.265 180.215 ;
        RECT 64.860 180.100 65.310 183.775 ;
        RECT 82.690 181.440 83.140 185.515 ;
        RECT 83.960 185.465 98.465 185.515 ;
        RECT 84.860 185.405 98.465 185.465 ;
        RECT 85.765 185.345 98.465 185.405 ;
        RECT 85.765 185.330 99.345 185.345 ;
        RECT 86.665 185.245 99.345 185.330 ;
        RECT 87.565 185.150 99.345 185.245 ;
        RECT 88.460 185.115 99.345 185.150 ;
        RECT 88.460 185.040 100.220 185.115 ;
        RECT 89.360 184.920 100.220 185.040 ;
        RECT 90.255 184.875 100.220 184.920 ;
        RECT 90.255 184.790 101.090 184.875 ;
        RECT 91.145 184.650 101.090 184.790 ;
        RECT 92.040 184.620 101.090 184.650 ;
        RECT 92.040 184.495 101.960 184.620 ;
        RECT 92.930 184.360 101.960 184.495 ;
        RECT 92.930 184.330 102.825 184.360 ;
        RECT 93.815 184.155 102.825 184.330 ;
        RECT 94.700 184.085 102.825 184.155 ;
        RECT 94.700 183.970 103.685 184.085 ;
        RECT 95.585 183.800 103.685 183.970 ;
        RECT 95.585 183.775 104.545 183.800 ;
        RECT 96.465 183.565 104.545 183.775 ;
        RECT 97.345 183.505 104.545 183.565 ;
        RECT 97.345 183.345 105.400 183.505 ;
        RECT 98.220 183.195 105.400 183.345 ;
        RECT 98.220 183.115 106.250 183.195 ;
        RECT 99.090 182.880 106.250 183.115 ;
        RECT 99.090 182.875 107.100 182.880 ;
        RECT 99.960 182.620 107.100 182.875 ;
        RECT 85.170 182.210 87.570 182.510 ;
        RECT 84.870 181.910 87.570 182.210 ;
        RECT 84.270 181.310 88.170 181.910 ;
        RECT 67.340 180.870 69.740 181.170 ;
        RECT 67.040 180.570 69.740 180.870 ;
        RECT 66.440 179.970 70.340 180.570 ;
        RECT 83.970 180.110 88.470 181.310 ;
        RECT 47.160 179.865 53.265 179.965 ;
        RECT 47.160 179.555 52.435 179.865 ;
        RECT 46.355 179.505 52.435 179.555 ;
        RECT 46.355 179.135 51.605 179.505 ;
        RECT 46.355 179.130 50.785 179.135 ;
        RECT 45.550 178.755 50.785 179.130 ;
        RECT 66.140 178.770 70.640 179.970 ;
        RECT 83.970 179.810 84.870 180.110 ;
        RECT 83.970 179.510 84.570 179.810 ;
        RECT 45.550 178.700 49.970 178.755 ;
        RECT 44.755 178.365 49.970 178.700 ;
        RECT 66.140 178.470 67.040 178.770 ;
        RECT 44.755 178.260 49.160 178.365 ;
        RECT 43.965 177.965 49.160 178.260 ;
        RECT 66.140 178.170 66.740 178.470 ;
        RECT 43.965 177.810 48.670 177.965 ;
        RECT 43.180 177.555 48.670 177.810 ;
        RECT 43.180 177.350 47.550 177.555 ;
        RECT 42.405 177.130 47.550 177.350 ;
        RECT 42.405 176.880 46.755 177.130 ;
        RECT 41.630 176.700 46.755 176.880 ;
        RECT 41.630 176.400 45.965 176.700 ;
        RECT 40.865 176.260 45.965 176.400 ;
        RECT 40.865 175.910 45.180 176.260 ;
        RECT 40.100 175.810 45.180 175.910 ;
        RECT 40.100 175.410 44.405 175.810 ;
        RECT 39.345 175.350 44.405 175.410 ;
        RECT 39.345 174.900 43.630 175.350 ;
        RECT 38.600 174.880 43.630 174.900 ;
        RECT 38.600 174.400 42.865 174.880 ;
        RECT 38.600 174.385 42.100 174.400 ;
        RECT 37.855 173.910 42.100 174.385 ;
        RECT 37.855 173.855 41.345 173.910 ;
        RECT 37.120 173.410 41.345 173.855 ;
        RECT 48.220 173.570 48.670 177.555 ;
        RECT 66.440 177.870 66.740 178.170 ;
        RECT 67.940 177.870 68.840 178.770 ;
        RECT 69.740 178.470 70.640 178.770 ;
        RECT 84.270 179.210 84.570 179.510 ;
        RECT 85.770 179.210 86.670 180.110 ;
        RECT 87.570 179.810 88.470 180.110 ;
        RECT 87.870 179.510 88.470 179.810 ;
        RECT 87.870 179.210 88.170 179.510 ;
        RECT 84.270 178.910 84.870 179.210 ;
        RECT 85.470 178.910 86.970 179.210 ;
        RECT 87.570 178.910 88.170 179.210 ;
        RECT 84.270 178.610 86.070 178.910 ;
        RECT 86.370 178.610 87.870 178.910 ;
        RECT 70.040 178.170 70.640 178.470 ;
        RECT 84.870 178.310 85.770 178.610 ;
        RECT 86.670 178.310 87.870 178.610 ;
        RECT 70.040 177.870 70.340 178.170 ;
        RECT 66.440 177.570 67.040 177.870 ;
        RECT 67.640 177.570 69.140 177.870 ;
        RECT 69.740 177.570 70.340 177.870 ;
        RECT 85.170 177.710 87.270 178.310 ;
        RECT 66.440 177.270 68.240 177.570 ;
        RECT 68.540 177.270 70.040 177.570 ;
        RECT 83.370 177.410 84.270 177.710 ;
        RECT 85.170 177.410 85.470 177.710 ;
        RECT 85.770 177.410 86.070 177.710 ;
        RECT 86.370 177.410 86.670 177.710 ;
        RECT 86.970 177.410 87.270 177.710 ;
        RECT 88.170 177.410 89.070 177.710 ;
        RECT 100.130 177.460 100.580 182.620 ;
        RECT 100.825 182.550 107.100 182.620 ;
        RECT 100.825 182.360 107.940 182.550 ;
        RECT 101.685 182.215 107.940 182.360 ;
        RECT 101.685 182.085 108.780 182.215 ;
        RECT 102.545 181.865 108.780 182.085 ;
        RECT 102.545 181.800 109.615 181.865 ;
        RECT 103.400 181.505 109.615 181.800 ;
        RECT 104.250 181.195 110.445 181.505 ;
        RECT 105.100 181.135 110.445 181.195 ;
        RECT 105.100 180.880 111.275 181.135 ;
        RECT 105.940 180.755 111.275 180.880 ;
        RECT 105.940 180.550 112.095 180.755 ;
        RECT 106.780 180.365 112.095 180.550 ;
        RECT 106.780 180.215 112.910 180.365 ;
        RECT 107.615 179.965 112.910 180.215 ;
        RECT 107.615 179.865 113.720 179.965 ;
        RECT 108.445 179.555 113.720 179.865 ;
        RECT 108.445 179.505 114.525 179.555 ;
        RECT 109.275 179.135 114.525 179.505 ;
        RECT 110.095 179.130 114.525 179.135 ;
        RECT 110.095 178.755 115.330 179.130 ;
        RECT 110.910 178.700 115.330 178.755 ;
        RECT 102.610 178.230 105.010 178.530 ;
        RECT 110.910 178.365 116.125 178.700 ;
        RECT 102.310 177.930 105.010 178.230 ;
        RECT 111.720 178.260 116.125 178.365 ;
        RECT 111.720 177.965 116.915 178.260 ;
        RECT 67.040 176.970 67.940 177.270 ;
        RECT 68.840 176.970 70.040 177.270 ;
        RECT 67.340 176.370 69.440 176.970 ;
        RECT 83.070 176.810 84.570 177.410 ;
        RECT 87.870 176.810 89.370 177.410 ;
        RECT 101.710 177.330 105.610 177.930 ;
        RECT 112.525 177.810 116.915 177.965 ;
        RECT 112.525 177.555 117.700 177.810 ;
        RECT 113.330 177.350 117.700 177.555 ;
        RECT 83.370 176.510 85.170 176.810 ;
        RECT 87.270 176.510 89.070 176.810 ;
        RECT 65.540 176.070 66.440 176.370 ;
        RECT 67.340 176.070 67.640 176.370 ;
        RECT 67.940 176.070 68.240 176.370 ;
        RECT 68.540 176.070 68.840 176.370 ;
        RECT 69.140 176.070 69.440 176.370 ;
        RECT 70.340 176.070 71.240 176.370 ;
        RECT 84.270 176.210 85.470 176.510 ;
        RECT 86.970 176.210 88.170 176.510 ;
        RECT 65.240 175.470 66.740 176.070 ;
        RECT 70.040 175.470 71.540 176.070 ;
        RECT 84.870 175.910 86.070 176.210 ;
        RECT 86.370 175.910 87.570 176.210 ;
        RECT 101.410 176.130 105.910 177.330 ;
        RECT 113.330 177.130 118.475 177.350 ;
        RECT 114.125 176.880 118.475 177.130 ;
        RECT 114.125 176.700 119.250 176.880 ;
        RECT 114.915 176.400 119.250 176.700 ;
        RECT 114.915 176.260 120.015 176.400 ;
        RECT 65.540 175.170 67.340 175.470 ;
        RECT 69.440 175.170 71.240 175.470 ;
        RECT 85.470 175.310 86.970 175.910 ;
        RECT 101.410 175.830 102.310 176.130 ;
        RECT 101.410 175.530 102.010 175.830 ;
        RECT 66.440 174.870 67.640 175.170 ;
        RECT 69.140 174.870 70.340 175.170 ;
        RECT 84.870 175.010 86.070 175.310 ;
        RECT 86.370 175.010 87.570 175.310 ;
        RECT 101.710 175.230 102.010 175.530 ;
        RECT 103.210 175.230 104.110 176.130 ;
        RECT 105.010 175.830 105.910 176.130 ;
        RECT 105.310 175.530 105.910 175.830 ;
        RECT 115.610 175.910 120.015 176.260 ;
        RECT 115.610 175.810 120.780 175.910 ;
        RECT 105.310 175.230 105.610 175.530 ;
        RECT 50.700 174.340 53.100 174.640 ;
        RECT 67.040 174.570 68.240 174.870 ;
        RECT 68.540 174.570 69.740 174.870 ;
        RECT 83.370 174.710 85.470 175.010 ;
        RECT 86.970 174.710 89.370 175.010 ;
        RECT 50.400 174.040 53.100 174.340 ;
        RECT 49.800 173.440 53.700 174.040 ;
        RECT 67.640 173.970 69.140 174.570 ;
        RECT 83.070 174.410 84.870 174.710 ;
        RECT 87.570 174.410 89.370 174.710 ;
        RECT 101.710 174.930 102.310 175.230 ;
        RECT 102.910 174.930 104.410 175.230 ;
        RECT 105.010 174.930 105.610 175.230 ;
        RECT 101.710 174.630 103.510 174.930 ;
        RECT 103.810 174.630 105.310 174.930 ;
        RECT 83.070 174.110 84.270 174.410 ;
        RECT 88.170 174.110 89.370 174.410 ;
        RECT 102.310 174.330 103.210 174.630 ;
        RECT 104.110 174.330 105.310 174.630 ;
        RECT 67.040 173.670 68.240 173.970 ;
        RECT 68.540 173.670 69.740 173.970 ;
        RECT 83.070 173.810 83.970 174.110 ;
        RECT 88.470 173.810 89.370 174.110 ;
        RECT 37.120 173.320 40.600 173.410 ;
        RECT 36.395 172.900 40.600 173.320 ;
        RECT 36.395 172.775 39.855 172.900 ;
        RECT 35.670 172.385 39.855 172.775 ;
        RECT 35.670 172.220 39.120 172.385 ;
        RECT 34.955 171.855 39.120 172.220 ;
        RECT 49.500 172.240 54.000 173.440 ;
        RECT 65.540 173.370 67.640 173.670 ;
        RECT 69.140 173.370 71.540 173.670 ;
        RECT 83.370 173.510 83.670 173.810 ;
        RECT 85.170 173.510 85.470 173.810 ;
        RECT 85.770 173.510 86.070 173.810 ;
        RECT 86.370 173.510 86.670 173.810 ;
        RECT 86.970 173.510 87.270 173.810 ;
        RECT 88.770 173.510 89.070 173.810 ;
        RECT 102.610 173.730 104.710 174.330 ;
        RECT 65.240 173.070 67.040 173.370 ;
        RECT 69.740 173.070 71.540 173.370 ;
        RECT 65.240 172.770 66.440 173.070 ;
        RECT 70.340 172.770 71.540 173.070 ;
        RECT 85.170 172.910 87.270 173.510 ;
        RECT 100.810 173.430 101.710 173.730 ;
        RECT 102.610 173.430 102.910 173.730 ;
        RECT 103.210 173.430 103.510 173.730 ;
        RECT 103.810 173.430 104.110 173.730 ;
        RECT 104.410 173.430 104.710 173.730 ;
        RECT 105.610 173.430 106.510 173.730 ;
        RECT 65.240 172.470 66.140 172.770 ;
        RECT 70.640 172.470 71.540 172.770 ;
        RECT 84.870 172.610 85.770 172.910 ;
        RECT 86.670 172.610 87.870 172.910 ;
        RECT 100.510 172.830 102.010 173.430 ;
        RECT 105.310 172.830 106.810 173.430 ;
        RECT 49.500 171.940 50.400 172.240 ;
        RECT 34.955 171.655 38.395 171.855 ;
        RECT 34.250 171.320 38.395 171.655 ;
        RECT 49.500 171.640 50.100 171.940 ;
        RECT 49.800 171.340 50.100 171.640 ;
        RECT 51.300 171.340 52.200 172.240 ;
        RECT 53.100 171.940 54.000 172.240 ;
        RECT 65.540 172.170 65.840 172.470 ;
        RECT 67.340 172.170 67.640 172.470 ;
        RECT 67.940 172.170 68.240 172.470 ;
        RECT 68.540 172.170 68.840 172.470 ;
        RECT 69.140 172.170 69.440 172.470 ;
        RECT 70.940 172.170 71.240 172.470 ;
        RECT 84.270 172.310 86.070 172.610 ;
        RECT 86.370 172.310 87.870 172.610 ;
        RECT 100.810 172.530 102.610 172.830 ;
        RECT 104.710 172.530 106.510 172.830 ;
        RECT 53.400 171.640 54.000 171.940 ;
        RECT 53.400 171.340 53.700 171.640 ;
        RECT 67.340 171.570 69.440 172.170 ;
        RECT 84.270 172.010 84.870 172.310 ;
        RECT 85.470 172.010 86.970 172.310 ;
        RECT 87.570 172.010 88.170 172.310 ;
        RECT 101.710 172.230 102.910 172.530 ;
        RECT 104.410 172.230 105.610 172.530 ;
        RECT 84.270 171.710 84.570 172.010 ;
        RECT 34.250 171.085 37.670 171.320 ;
        RECT 33.550 170.775 37.670 171.085 ;
        RECT 49.800 171.040 50.400 171.340 ;
        RECT 51.000 171.040 52.500 171.340 ;
        RECT 53.100 171.040 53.700 171.340 ;
        RECT 67.040 171.270 67.940 171.570 ;
        RECT 68.840 171.270 70.040 171.570 ;
        RECT 33.550 170.505 36.955 170.775 ;
        RECT 49.800 170.740 51.600 171.040 ;
        RECT 51.900 170.740 53.400 171.040 ;
        RECT 32.855 170.220 36.955 170.505 ;
        RECT 50.400 170.440 51.300 170.740 ;
        RECT 52.200 170.440 53.400 170.740 ;
        RECT 66.440 170.970 68.240 171.270 ;
        RECT 68.540 170.970 70.040 171.270 ;
        RECT 83.970 171.410 84.570 171.710 ;
        RECT 83.970 171.110 84.870 171.410 ;
        RECT 85.770 171.110 86.670 172.010 ;
        RECT 87.870 171.710 88.170 172.010 ;
        RECT 102.310 171.930 103.510 172.230 ;
        RECT 103.810 171.930 105.010 172.230 ;
        RECT 87.870 171.410 88.470 171.710 ;
        RECT 87.570 171.110 88.470 171.410 ;
        RECT 102.910 171.330 104.410 171.930 ;
        RECT 66.440 170.670 67.040 170.970 ;
        RECT 67.640 170.670 69.140 170.970 ;
        RECT 69.740 170.670 70.340 170.970 ;
        RECT 32.855 169.915 36.250 170.220 ;
        RECT 32.170 169.655 36.250 169.915 ;
        RECT 50.700 169.840 52.800 170.440 ;
        RECT 66.440 170.370 66.740 170.670 ;
        RECT 66.140 170.070 66.740 170.370 ;
        RECT 32.170 169.315 35.550 169.655 ;
        RECT 48.900 169.540 49.800 169.840 ;
        RECT 50.700 169.540 51.000 169.840 ;
        RECT 51.300 169.540 51.600 169.840 ;
        RECT 51.900 169.540 52.200 169.840 ;
        RECT 52.500 169.540 52.800 169.840 ;
        RECT 53.700 169.540 54.600 169.840 ;
        RECT 66.140 169.770 67.040 170.070 ;
        RECT 67.940 169.770 68.840 170.670 ;
        RECT 70.040 170.370 70.340 170.670 ;
        RECT 70.040 170.070 70.640 170.370 ;
        RECT 69.740 169.770 70.640 170.070 ;
        RECT 83.970 169.910 88.470 171.110 ;
        RECT 102.310 171.030 103.510 171.330 ;
        RECT 103.810 171.030 105.010 171.330 ;
        RECT 100.810 170.730 102.910 171.030 ;
        RECT 104.410 170.730 106.810 171.030 ;
        RECT 100.510 170.430 102.310 170.730 ;
        RECT 105.010 170.430 106.810 170.730 ;
        RECT 100.510 170.130 101.710 170.430 ;
        RECT 105.610 170.130 106.810 170.430 ;
        RECT 31.490 169.085 35.550 169.315 ;
        RECT 31.490 168.710 34.855 169.085 ;
        RECT 48.600 168.940 50.100 169.540 ;
        RECT 53.400 168.940 54.900 169.540 ;
        RECT 30.820 168.505 34.855 168.710 ;
        RECT 48.900 168.640 50.700 168.940 ;
        RECT 52.800 168.640 54.600 168.940 ;
        RECT 30.820 168.095 34.170 168.505 ;
        RECT 49.800 168.340 51.000 168.640 ;
        RECT 52.500 168.340 53.700 168.640 ;
        RECT 66.140 168.570 70.640 169.770 ;
        RECT 30.155 167.915 34.170 168.095 ;
        RECT 50.400 168.040 51.600 168.340 ;
        RECT 51.900 168.040 53.100 168.340 ;
        RECT 30.155 167.645 33.490 167.915 ;
        RECT 30.155 167.470 34.680 167.645 ;
        RECT 29.500 167.195 34.680 167.470 ;
        RECT 51.000 167.440 52.500 168.040 ;
        RECT 29.500 166.840 32.820 167.195 ;
        RECT 28.850 166.710 32.820 166.840 ;
        RECT 28.850 166.200 32.155 166.710 ;
        RECT 28.210 166.095 32.155 166.200 ;
        RECT 28.210 165.550 31.500 166.095 ;
        RECT 27.580 165.470 31.500 165.550 ;
        RECT 27.580 164.895 30.850 165.470 ;
        RECT 26.955 164.840 30.850 164.895 ;
        RECT 26.955 164.230 30.210 164.840 ;
        RECT 26.340 164.200 30.210 164.230 ;
        RECT 26.340 163.560 29.580 164.200 ;
        RECT 25.735 163.550 29.580 163.560 ;
        RECT 25.735 162.895 28.955 163.550 ;
        RECT 25.735 162.880 28.340 162.895 ;
        RECT 25.135 162.230 28.340 162.880 ;
        RECT 34.230 162.420 34.680 167.195 ;
        RECT 50.400 167.140 51.600 167.440 ;
        RECT 51.900 167.140 53.100 167.440 ;
        RECT 48.900 166.840 51.000 167.140 ;
        RECT 52.500 166.840 54.900 167.140 ;
        RECT 48.600 166.540 50.400 166.840 ;
        RECT 53.100 166.540 54.900 166.840 ;
        RECT 48.600 166.240 49.800 166.540 ;
        RECT 53.700 166.240 54.900 166.540 ;
        RECT 48.600 165.940 49.500 166.240 ;
        RECT 54.000 165.940 54.900 166.240 ;
        RECT 64.860 166.980 65.420 168.370 ;
        RECT 66.440 167.970 70.340 168.570 ;
        RECT 82.690 168.320 83.250 169.710 ;
        RECT 84.270 169.310 88.170 169.910 ;
        RECT 100.510 169.830 101.410 170.130 ;
        RECT 105.910 169.830 106.810 170.130 ;
        RECT 100.810 169.530 101.110 169.830 ;
        RECT 102.610 169.530 102.910 169.830 ;
        RECT 103.210 169.530 103.510 169.830 ;
        RECT 103.810 169.530 104.110 169.830 ;
        RECT 104.410 169.530 104.710 169.830 ;
        RECT 106.210 169.530 106.510 169.830 ;
        RECT 84.870 169.010 87.570 169.310 ;
        RECT 85.170 168.710 87.570 169.010 ;
        RECT 102.610 168.930 104.710 169.530 ;
        RECT 102.310 168.630 103.210 168.930 ;
        RECT 104.110 168.630 105.310 168.930 ;
        RECT 101.710 168.330 103.510 168.630 ;
        RECT 103.810 168.330 105.310 168.630 ;
        RECT 115.610 168.510 116.060 175.810 ;
        RECT 116.475 175.410 120.780 175.810 ;
        RECT 116.475 175.350 121.535 175.410 ;
        RECT 117.250 174.900 121.535 175.350 ;
        RECT 117.250 174.880 122.280 174.900 ;
        RECT 118.015 174.400 122.280 174.880 ;
        RECT 118.780 174.385 122.280 174.400 ;
        RECT 118.780 173.910 123.025 174.385 ;
        RECT 119.535 173.855 123.025 173.910 ;
        RECT 119.535 173.410 123.760 173.855 ;
        RECT 120.280 173.320 123.760 173.410 ;
        RECT 120.280 172.900 124.485 173.320 ;
        RECT 121.025 172.775 124.485 172.900 ;
        RECT 121.025 172.385 125.210 172.775 ;
        RECT 121.760 172.220 125.210 172.385 ;
        RECT 121.760 171.855 125.925 172.220 ;
        RECT 122.485 171.655 125.925 171.855 ;
        RECT 122.485 171.320 126.630 171.655 ;
        RECT 123.210 171.085 126.630 171.320 ;
        RECT 123.210 170.775 127.330 171.085 ;
        RECT 123.925 170.505 127.330 170.775 ;
        RECT 123.925 170.220 128.025 170.505 ;
        RECT 124.630 169.915 128.025 170.220 ;
        RECT 124.630 169.655 128.710 169.915 ;
        RECT 118.090 169.280 120.490 169.580 ;
        RECT 117.790 168.980 120.490 169.280 ;
        RECT 125.330 169.315 128.710 169.655 ;
        RECT 125.330 169.085 129.390 169.315 ;
        RECT 117.190 168.380 121.090 168.980 ;
        RECT 126.025 168.710 129.390 169.085 ;
        RECT 126.025 168.505 130.060 168.710 ;
        RECT 67.040 167.670 69.740 167.970 ;
        RECT 67.340 167.370 69.740 167.670 ;
        RECT 48.900 165.640 49.200 165.940 ;
        RECT 50.700 165.640 51.000 165.940 ;
        RECT 51.300 165.640 51.600 165.940 ;
        RECT 51.900 165.640 52.200 165.940 ;
        RECT 52.500 165.640 52.800 165.940 ;
        RECT 54.300 165.640 54.600 165.940 ;
        RECT 50.700 165.040 52.800 165.640 ;
        RECT 50.400 164.740 51.300 165.040 ;
        RECT 52.200 164.740 53.400 165.040 ;
        RECT 49.800 164.440 51.600 164.740 ;
        RECT 51.900 164.440 53.400 164.740 ;
        RECT 49.800 164.140 50.400 164.440 ;
        RECT 51.000 164.140 52.500 164.440 ;
        RECT 53.100 164.140 53.700 164.440 ;
        RECT 49.800 163.840 50.100 164.140 ;
        RECT 49.500 163.540 50.100 163.840 ;
        RECT 36.710 163.190 39.110 163.490 ;
        RECT 36.410 162.890 39.110 163.190 ;
        RECT 49.500 163.240 50.400 163.540 ;
        RECT 51.300 163.240 52.200 164.140 ;
        RECT 53.400 163.840 53.700 164.140 ;
        RECT 53.400 163.540 54.000 163.840 ;
        RECT 53.100 163.240 54.000 163.540 ;
        RECT 35.810 162.290 39.710 162.890 ;
        RECT 25.135 162.195 27.735 162.230 ;
        RECT 24.545 161.560 27.735 162.195 ;
        RECT 24.545 161.500 27.135 161.560 ;
        RECT 23.965 160.880 27.135 161.500 ;
        RECT 35.510 161.090 40.010 162.290 ;
        RECT 49.500 162.040 54.000 163.240 ;
        RECT 64.860 162.465 65.310 166.980 ;
        RECT 79.445 164.600 81.440 164.610 ;
        RECT 78.585 164.580 82.295 164.600 ;
        RECT 82.690 164.580 83.140 168.320 ;
        RECT 101.710 168.030 102.310 168.330 ;
        RECT 102.910 168.030 104.410 168.330 ;
        RECT 105.010 168.030 105.610 168.330 ;
        RECT 101.710 167.730 102.010 168.030 ;
        RECT 101.410 167.430 102.010 167.730 ;
        RECT 101.410 167.130 102.310 167.430 ;
        RECT 103.210 167.130 104.110 168.030 ;
        RECT 105.310 167.730 105.610 168.030 ;
        RECT 105.310 167.430 105.910 167.730 ;
        RECT 105.010 167.130 105.910 167.430 ;
        RECT 101.410 165.930 105.910 167.130 ;
        RECT 116.890 167.180 121.390 168.380 ;
        RECT 126.710 168.095 130.060 168.505 ;
        RECT 126.710 167.915 130.725 168.095 ;
        RECT 127.390 167.470 130.725 167.915 ;
        RECT 127.390 167.315 131.380 167.470 ;
        RECT 116.890 166.880 117.790 167.180 ;
        RECT 116.890 166.580 117.490 166.880 ;
        RECT 117.190 166.280 117.490 166.580 ;
        RECT 118.690 166.280 119.590 167.180 ;
        RECT 120.490 166.880 121.390 167.180 ;
        RECT 120.790 166.580 121.390 166.880 ;
        RECT 128.060 166.840 131.380 167.315 ;
        RECT 128.060 166.710 132.030 166.840 ;
        RECT 120.790 166.280 121.090 166.580 ;
        RECT 117.190 165.980 117.790 166.280 ;
        RECT 118.390 165.980 119.890 166.280 ;
        RECT 120.490 165.980 121.090 166.280 ;
        RECT 128.725 166.200 132.030 166.710 ;
        RECT 128.725 166.095 132.670 166.200 ;
        RECT 77.730 164.540 83.150 164.580 ;
        RECT 76.880 164.490 84.000 164.540 ;
        RECT 76.025 164.420 84.855 164.490 ;
        RECT 75.170 164.340 85.710 164.420 ;
        RECT 100.130 164.340 100.690 165.730 ;
        RECT 101.710 165.330 105.610 165.930 ;
        RECT 117.190 165.680 118.990 165.980 ;
        RECT 119.290 165.680 120.790 165.980 ;
        RECT 117.790 165.380 118.690 165.680 ;
        RECT 119.590 165.380 120.790 165.680 ;
        RECT 129.380 165.550 132.670 166.095 ;
        RECT 129.380 165.470 133.300 165.550 ;
        RECT 102.310 165.030 105.010 165.330 ;
        RECT 102.610 164.730 105.010 165.030 ;
        RECT 118.090 164.780 120.190 165.380 ;
        RECT 130.030 164.895 133.300 165.470 ;
        RECT 130.030 164.840 133.925 164.895 ;
        RECT 116.290 164.480 117.190 164.780 ;
        RECT 118.090 164.480 118.390 164.780 ;
        RECT 118.690 164.480 118.990 164.780 ;
        RECT 119.290 164.480 119.590 164.780 ;
        RECT 119.890 164.480 120.190 164.780 ;
        RECT 121.090 164.480 121.990 164.780 ;
        RECT 74.320 164.240 86.560 164.340 ;
        RECT 73.470 164.130 87.410 164.240 ;
        RECT 72.625 164.005 88.255 164.130 ;
        RECT 71.775 163.865 89.105 164.005 ;
        RECT 70.935 163.705 89.945 163.865 ;
        RECT 70.095 163.535 90.785 163.705 ;
        RECT 69.255 163.350 91.625 163.535 ;
        RECT 68.420 163.150 92.460 163.350 ;
        RECT 67.590 162.940 93.290 163.150 ;
        RECT 66.760 162.710 94.120 162.940 ;
        RECT 65.935 162.600 94.945 162.710 ;
        RECT 65.935 162.580 79.730 162.600 ;
        RECT 81.150 162.580 94.945 162.600 ;
        RECT 65.935 162.540 78.880 162.580 ;
        RECT 82.000 162.540 94.945 162.580 ;
        RECT 65.935 162.490 78.025 162.540 ;
        RECT 82.855 162.490 94.945 162.540 ;
        RECT 65.935 162.465 77.170 162.490 ;
        RECT 64.860 162.420 77.170 162.465 ;
        RECT 83.710 162.465 94.945 162.490 ;
        RECT 83.710 162.420 95.765 162.465 ;
        RECT 64.860 162.340 76.320 162.420 ;
        RECT 84.560 162.340 95.765 162.420 ;
        RECT 64.860 162.240 75.470 162.340 ;
        RECT 85.410 162.240 95.765 162.340 ;
        RECT 64.860 162.210 74.625 162.240 ;
        RECT 64.300 162.130 74.625 162.210 ;
        RECT 86.255 162.210 95.765 162.240 ;
        RECT 86.255 162.130 96.580 162.210 ;
        RECT 23.965 160.800 26.545 160.880 ;
        RECT 23.395 160.195 26.545 160.800 ;
        RECT 35.510 160.790 36.410 161.090 ;
        RECT 35.510 160.490 36.110 160.790 ;
        RECT 23.395 160.095 25.965 160.195 ;
        RECT 22.830 159.500 25.965 160.095 ;
        RECT 35.810 160.190 36.110 160.490 ;
        RECT 37.310 160.190 38.210 161.090 ;
        RECT 39.110 160.790 40.010 161.090 ;
        RECT 39.410 160.490 40.010 160.790 ;
        RECT 39.410 160.190 39.710 160.490 ;
        RECT 35.810 159.890 36.410 160.190 ;
        RECT 37.010 159.890 38.510 160.190 ;
        RECT 39.110 159.890 39.710 160.190 ;
        RECT 48.220 160.450 48.780 161.840 ;
        RECT 49.800 161.440 53.700 162.040 ;
        RECT 64.300 162.005 73.775 162.130 ;
        RECT 87.105 162.005 96.580 162.130 ;
        RECT 64.300 161.940 72.935 162.005 ;
        RECT 63.490 161.865 72.935 161.940 ;
        RECT 87.945 161.940 96.580 162.005 ;
        RECT 87.945 161.865 97.390 161.940 ;
        RECT 63.490 161.705 72.095 161.865 ;
        RECT 88.785 161.705 97.390 161.865 ;
        RECT 63.490 161.650 71.255 161.705 ;
        RECT 62.685 161.535 71.255 161.650 ;
        RECT 89.625 161.650 97.390 161.705 ;
        RECT 89.625 161.535 98.195 161.650 ;
        RECT 50.400 161.140 53.100 161.440 ;
        RECT 62.685 161.355 70.420 161.535 ;
        RECT 50.700 160.840 53.100 161.140 ;
        RECT 61.880 161.350 70.420 161.355 ;
        RECT 90.460 161.355 98.195 161.535 ;
        RECT 90.460 161.350 99.000 161.355 ;
        RECT 61.880 161.150 69.590 161.350 ;
        RECT 91.290 161.150 99.000 161.350 ;
        RECT 61.880 161.040 68.760 161.150 ;
        RECT 61.085 160.940 68.760 161.040 ;
        RECT 92.120 161.040 99.000 161.150 ;
        RECT 92.120 160.940 99.795 161.040 ;
        RECT 61.085 160.710 67.935 160.940 ;
        RECT 92.945 160.710 99.795 160.940 ;
        RECT 100.130 160.710 100.580 164.340 ;
        RECT 115.990 163.880 117.490 164.480 ;
        RECT 120.790 163.880 122.290 164.480 ;
        RECT 130.670 164.230 133.925 164.840 ;
        RECT 130.670 164.200 134.540 164.230 ;
        RECT 116.290 163.580 118.090 163.880 ;
        RECT 120.190 163.580 121.990 163.880 ;
        RECT 117.190 163.280 118.390 163.580 ;
        RECT 119.890 163.280 121.090 163.580 ;
        RECT 131.300 163.560 134.540 164.200 ;
        RECT 131.300 163.550 135.145 163.560 ;
        RECT 117.790 162.980 118.990 163.280 ;
        RECT 119.290 162.980 120.490 163.280 ;
        RECT 118.390 162.380 119.890 162.980 ;
        RECT 131.925 162.895 135.145 163.550 ;
        RECT 132.540 162.880 135.145 162.895 ;
        RECT 117.790 162.080 118.990 162.380 ;
        RECT 119.290 162.080 120.490 162.380 ;
        RECT 132.540 162.230 135.745 162.880 ;
        RECT 133.145 162.195 135.745 162.230 ;
        RECT 116.290 161.780 118.390 162.080 ;
        RECT 119.890 161.780 122.290 162.080 ;
        RECT 115.990 161.480 117.790 161.780 ;
        RECT 120.490 161.480 122.290 161.780 ;
        RECT 133.145 161.560 136.335 162.195 ;
        RECT 115.990 161.180 117.190 161.480 ;
        RECT 121.090 161.180 122.290 161.480 ;
        RECT 115.990 160.880 116.890 161.180 ;
        RECT 121.390 160.880 122.290 161.180 ;
        RECT 133.745 161.500 136.335 161.560 ;
        RECT 133.745 160.880 136.915 161.500 ;
        RECT 60.295 160.465 67.115 160.710 ;
        RECT 93.765 160.465 100.585 160.710 ;
        RECT 116.290 160.580 116.590 160.880 ;
        RECT 118.090 160.580 118.390 160.880 ;
        RECT 118.690 160.580 118.990 160.880 ;
        RECT 119.290 160.580 119.590 160.880 ;
        RECT 119.890 160.580 120.190 160.880 ;
        RECT 121.690 160.580 121.990 160.880 ;
        RECT 134.335 160.800 136.915 160.880 ;
        RECT 35.810 159.590 37.610 159.890 ;
        RECT 37.910 159.590 39.410 159.890 ;
        RECT 22.830 159.380 25.395 159.500 ;
        RECT 22.275 158.800 25.395 159.380 ;
        RECT 36.410 159.290 37.310 159.590 ;
        RECT 38.210 159.290 39.410 159.590 ;
        RECT 22.275 158.655 24.830 158.800 ;
        RECT 36.710 158.690 38.810 159.290 ;
        RECT 21.730 158.095 24.830 158.655 ;
        RECT 34.910 158.390 35.810 158.690 ;
        RECT 36.710 158.390 37.010 158.690 ;
        RECT 37.310 158.390 37.610 158.690 ;
        RECT 37.910 158.390 38.210 158.690 ;
        RECT 38.510 158.390 38.810 158.690 ;
        RECT 39.710 158.390 40.610 158.690 ;
        RECT 21.730 157.930 24.275 158.095 ;
        RECT 21.195 157.380 24.275 157.930 ;
        RECT 34.610 157.790 36.110 158.390 ;
        RECT 39.410 157.790 40.910 158.390 ;
        RECT 34.910 157.490 36.710 157.790 ;
        RECT 38.810 157.490 40.610 157.790 ;
        RECT 21.195 157.195 23.730 157.380 ;
        RECT 20.665 156.655 23.730 157.195 ;
        RECT 35.810 157.190 37.010 157.490 ;
        RECT 38.510 157.190 39.710 157.490 ;
        RECT 36.410 156.890 37.610 157.190 ;
        RECT 37.910 156.890 39.110 157.190 ;
        RECT 20.665 156.450 23.195 156.655 ;
        RECT 20.150 155.930 23.195 156.450 ;
        RECT 37.010 156.290 38.510 156.890 ;
        RECT 36.410 155.990 37.610 156.290 ;
        RECT 37.910 155.990 39.110 156.290 ;
        RECT 20.150 155.705 22.665 155.930 ;
        RECT 19.640 155.195 22.665 155.705 ;
        RECT 34.910 155.690 37.010 155.990 ;
        RECT 38.510 155.690 40.910 155.990 ;
        RECT 34.610 155.390 36.410 155.690 ;
        RECT 39.110 155.390 40.910 155.690 ;
        RECT 19.640 154.950 22.150 155.195 ;
        RECT 19.140 154.450 22.150 154.950 ;
        RECT 34.610 155.090 35.810 155.390 ;
        RECT 39.710 155.090 40.910 155.390 ;
        RECT 34.610 154.790 35.510 155.090 ;
        RECT 40.010 154.790 40.910 155.090 ;
        RECT 34.910 154.490 35.210 154.790 ;
        RECT 36.710 154.490 37.010 154.790 ;
        RECT 37.310 154.490 37.610 154.790 ;
        RECT 37.910 154.490 38.210 154.790 ;
        RECT 38.510 154.490 38.810 154.790 ;
        RECT 40.310 154.490 40.610 154.790 ;
        RECT 19.140 154.185 21.640 154.450 ;
        RECT 18.650 153.705 21.640 154.185 ;
        RECT 36.710 153.890 38.810 154.490 ;
        RECT 18.650 153.420 21.140 153.705 ;
        RECT 36.410 153.590 37.310 153.890 ;
        RECT 38.210 153.590 39.410 153.890 ;
        RECT 18.170 152.950 21.140 153.420 ;
        RECT 35.810 153.290 37.610 153.590 ;
        RECT 37.910 153.290 39.410 153.590 ;
        RECT 48.220 153.690 48.670 160.450 ;
        RECT 60.295 160.370 66.300 160.465 ;
        RECT 59.510 160.210 66.300 160.370 ;
        RECT 94.580 160.370 100.585 160.465 ;
        RECT 94.580 160.210 101.370 160.370 ;
        RECT 59.510 160.015 65.490 160.210 ;
        RECT 58.735 159.940 65.490 160.015 ;
        RECT 95.390 160.015 101.370 160.210 ;
        RECT 95.390 159.940 102.145 160.015 ;
        RECT 118.090 159.980 120.190 160.580 ;
        RECT 134.335 160.195 137.485 160.800 ;
        RECT 134.915 160.095 137.485 160.195 ;
        RECT 58.735 159.650 64.685 159.940 ;
        RECT 96.195 159.650 102.145 159.940 ;
        RECT 117.790 159.680 118.690 159.980 ;
        RECT 119.590 159.680 120.790 159.980 ;
        RECT 57.960 159.355 63.880 159.650 ;
        RECT 97.000 159.355 102.920 159.650 ;
        RECT 57.960 159.265 63.085 159.355 ;
        RECT 57.195 159.040 63.085 159.265 ;
        RECT 97.795 159.265 102.920 159.355 ;
        RECT 117.190 159.380 118.990 159.680 ;
        RECT 119.290 159.380 120.790 159.680 ;
        RECT 134.915 159.500 138.050 160.095 ;
        RECT 135.485 159.380 138.050 159.500 ;
        RECT 97.795 159.040 103.685 159.265 ;
        RECT 57.195 158.870 62.295 159.040 ;
        RECT 56.440 158.710 62.295 158.870 ;
        RECT 98.585 158.870 103.685 159.040 ;
        RECT 117.190 159.080 117.790 159.380 ;
        RECT 118.390 159.080 119.890 159.380 ;
        RECT 120.490 159.080 121.090 159.380 ;
        RECT 98.585 158.710 104.440 158.870 ;
        RECT 117.190 158.780 117.490 159.080 ;
        RECT 56.440 158.465 61.510 158.710 ;
        RECT 55.685 158.370 61.510 158.465 ;
        RECT 99.370 158.465 104.440 158.710 ;
        RECT 116.890 158.480 117.490 158.780 ;
        RECT 99.370 158.370 105.195 158.465 ;
        RECT 55.685 158.045 60.735 158.370 ;
        RECT 54.945 158.015 60.735 158.045 ;
        RECT 100.145 158.045 105.195 158.370 ;
        RECT 116.890 158.180 117.790 158.480 ;
        RECT 118.690 158.180 119.590 159.080 ;
        RECT 120.790 158.780 121.090 159.080 ;
        RECT 135.485 158.800 138.605 159.380 ;
        RECT 120.790 158.480 121.390 158.780 ;
        RECT 120.490 158.180 121.390 158.480 ;
        RECT 100.145 158.015 105.940 158.045 ;
        RECT 54.945 157.650 59.960 158.015 ;
        RECT 100.920 157.650 105.940 158.015 ;
        RECT 54.945 157.610 59.195 157.650 ;
        RECT 54.205 157.265 59.195 157.610 ;
        RECT 101.685 157.610 105.940 157.650 ;
        RECT 101.685 157.265 106.675 157.610 ;
        RECT 54.205 157.160 58.440 157.265 ;
        RECT 53.475 156.870 58.440 157.160 ;
        RECT 102.440 157.160 106.675 157.265 ;
        RECT 102.440 156.870 107.405 157.160 ;
        RECT 116.890 156.980 121.390 158.180 ;
        RECT 136.050 158.655 138.605 158.800 ;
        RECT 136.050 158.095 139.150 158.655 ;
        RECT 136.605 157.930 139.150 158.095 ;
        RECT 136.605 157.765 139.685 157.930 ;
        RECT 127.780 157.315 139.685 157.765 ;
        RECT 53.475 156.700 57.685 156.870 ;
        RECT 52.755 156.465 57.685 156.700 ;
        RECT 103.195 156.700 107.405 156.870 ;
        RECT 103.195 156.465 108.125 156.700 ;
        RECT 52.755 156.230 56.945 156.465 ;
        RECT 52.040 156.045 56.945 156.230 ;
        RECT 103.940 156.230 108.125 156.465 ;
        RECT 103.940 156.045 108.840 156.230 ;
        RECT 52.040 155.745 56.205 156.045 ;
        RECT 51.335 155.610 56.205 155.745 ;
        RECT 104.675 155.745 108.840 156.045 ;
        RECT 104.675 155.610 109.545 155.745 ;
        RECT 51.335 155.250 55.475 155.610 ;
        RECT 50.640 155.160 55.475 155.250 ;
        RECT 105.405 155.250 109.545 155.610 ;
        RECT 115.610 155.390 116.170 156.780 ;
        RECT 117.190 156.380 121.090 156.980 ;
        RECT 117.790 156.080 120.490 156.380 ;
        RECT 118.090 155.780 120.490 156.080 ;
        RECT 127.780 155.400 128.230 157.315 ;
        RECT 137.150 157.195 139.685 157.315 ;
        RECT 137.150 156.655 140.215 157.195 ;
        RECT 130.260 156.170 132.660 156.470 ;
        RECT 129.960 155.870 132.660 156.170 ;
        RECT 137.685 156.450 140.215 156.655 ;
        RECT 137.685 155.930 140.730 156.450 ;
        RECT 105.405 155.160 110.240 155.250 ;
        RECT 50.640 154.740 54.755 155.160 ;
        RECT 49.955 154.700 54.755 154.740 ;
        RECT 49.955 154.230 54.040 154.700 ;
        RECT 49.955 154.220 53.335 154.230 ;
        RECT 49.275 153.745 53.335 154.220 ;
        RECT 49.275 153.690 52.640 153.745 ;
        RECT 35.810 152.990 36.410 153.290 ;
        RECT 37.010 152.990 38.510 153.290 ;
        RECT 39.110 152.990 39.710 153.290 ;
        RECT 48.220 153.250 52.640 153.690 ;
        RECT 48.220 153.145 51.955 153.250 ;
        RECT 18.170 152.645 20.650 152.950 ;
        RECT 35.810 152.690 36.110 152.990 ;
        RECT 17.700 152.185 20.650 152.645 ;
        RECT 35.510 152.390 36.110 152.690 ;
        RECT 17.700 151.870 20.170 152.185 ;
        RECT 17.240 151.420 20.170 151.870 ;
        RECT 35.510 152.090 36.410 152.390 ;
        RECT 37.310 152.090 38.210 152.990 ;
        RECT 39.410 152.690 39.710 152.990 ;
        RECT 47.945 152.740 51.955 153.145 ;
        RECT 39.410 152.390 40.010 152.690 ;
        RECT 47.945 152.590 51.275 152.740 ;
        RECT 39.110 152.090 40.010 152.390 ;
        RECT 17.240 151.085 19.700 151.420 ;
        RECT 16.790 150.645 19.700 151.085 ;
        RECT 35.510 150.890 40.010 152.090 ;
        RECT 47.295 152.220 51.275 152.590 ;
        RECT 47.295 152.020 50.605 152.220 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 106.125 154.740 110.240 155.160 ;
        RECT 106.125 154.700 110.925 154.740 ;
        RECT 106.840 154.230 110.925 154.700 ;
        RECT 107.545 154.220 110.925 154.230 ;
        RECT 107.545 153.745 111.605 154.220 ;
        RECT 108.240 153.690 111.605 153.745 ;
        RECT 108.240 153.250 112.275 153.690 ;
        RECT 108.925 153.145 112.275 153.250 ;
        RECT 108.925 152.740 112.935 153.145 ;
        RECT 109.605 152.590 112.935 152.740 ;
        RECT 109.605 152.220 113.585 152.590 ;
        RECT 115.610 152.255 116.060 155.390 ;
        RECT 129.360 155.270 133.260 155.870 ;
        RECT 138.215 155.705 140.730 155.930 ;
        RECT 129.060 154.070 133.560 155.270 ;
        RECT 138.215 155.195 141.240 155.705 ;
        RECT 138.730 154.950 141.240 155.195 ;
        RECT 138.730 154.450 141.740 154.950 ;
        RECT 129.060 153.770 129.960 154.070 ;
        RECT 129.060 153.470 129.660 153.770 ;
        RECT 129.360 153.170 129.660 153.470 ;
        RECT 130.860 153.170 131.760 154.070 ;
        RECT 132.660 153.770 133.560 154.070 ;
        RECT 132.960 153.470 133.560 153.770 ;
        RECT 139.240 154.185 141.740 154.450 ;
        RECT 139.240 153.705 142.230 154.185 ;
        RECT 132.960 153.170 133.260 153.470 ;
        RECT 129.360 152.870 129.960 153.170 ;
        RECT 130.560 152.870 132.060 153.170 ;
        RECT 132.660 152.870 133.260 153.170 ;
        RECT 139.740 153.420 142.230 153.705 ;
        RECT 139.740 152.950 142.710 153.420 ;
        RECT 129.360 152.570 131.160 152.870 ;
        RECT 131.460 152.570 132.960 152.870 ;
        RECT 129.960 152.270 130.860 152.570 ;
        RECT 131.760 152.270 132.960 152.570 ;
        RECT 140.230 152.645 142.710 152.950 ;
        RECT 46.655 151.690 50.605 152.020 ;
        RECT 46.655 151.445 49.945 151.690 ;
        RECT 46.025 151.145 49.945 151.445 ;
        RECT 16.790 150.295 19.240 150.645 ;
        RECT 16.350 149.870 19.240 150.295 ;
        RECT 16.350 149.640 18.790 149.870 ;
        RECT 16.350 149.500 24.610 149.640 ;
        RECT 15.920 149.190 24.610 149.500 ;
        RECT 15.920 149.085 18.790 149.190 ;
        RECT 15.920 148.695 18.350 149.085 ;
        RECT 15.495 148.295 18.350 148.695 ;
        RECT 15.495 147.890 17.920 148.295 ;
        RECT 15.085 147.500 17.920 147.890 ;
        RECT 24.160 147.640 24.610 149.190 ;
        RECT 34.230 149.300 34.790 150.690 ;
        RECT 35.810 150.290 39.710 150.890 ;
        RECT 46.025 150.855 49.295 151.145 ;
        RECT 45.405 150.590 49.295 150.855 ;
        RECT 36.410 149.990 39.110 150.290 ;
        RECT 45.405 150.255 48.655 150.590 ;
        RECT 36.710 149.690 39.110 149.990 ;
        RECT 44.795 150.020 48.655 150.255 ;
        RECT 44.795 149.645 48.025 150.020 ;
        RECT 44.195 149.445 48.025 149.645 ;
        RECT 68.170 149.600 91.570 152.200 ;
        RECT 110.275 152.020 113.585 152.220 ;
        RECT 110.275 151.690 114.225 152.020 ;
        RECT 110.935 151.445 114.225 151.690 ;
        RECT 110.935 151.145 114.855 151.445 ;
        RECT 111.585 150.855 114.855 151.145 ;
        RECT 115.605 150.855 116.065 152.255 ;
        RECT 130.260 151.670 132.360 152.270 ;
        RECT 140.230 152.185 143.180 152.645 ;
        RECT 140.710 151.870 143.180 152.185 ;
        RECT 128.460 151.370 129.360 151.670 ;
        RECT 130.260 151.370 130.560 151.670 ;
        RECT 130.860 151.370 131.160 151.670 ;
        RECT 131.460 151.370 131.760 151.670 ;
        RECT 132.060 151.370 132.360 151.670 ;
        RECT 133.260 151.370 134.160 151.670 ;
        RECT 140.710 151.420 143.640 151.870 ;
        RECT 111.585 150.590 116.065 150.855 ;
        RECT 128.160 150.770 129.660 151.370 ;
        RECT 132.960 150.770 134.460 151.370 ;
        RECT 141.180 151.085 143.640 151.420 ;
        RECT 112.225 150.255 116.065 150.590 ;
        RECT 128.460 150.470 130.260 150.770 ;
        RECT 132.360 150.470 134.160 150.770 ;
        RECT 141.180 150.645 144.090 151.085 ;
        RECT 112.225 150.020 116.085 150.255 ;
        RECT 129.360 150.170 130.560 150.470 ;
        RECT 132.060 150.170 133.260 150.470 ;
        RECT 141.640 150.295 144.090 150.645 ;
        RECT 112.855 149.645 116.085 150.020 ;
        RECT 129.960 149.870 131.160 150.170 ;
        RECT 131.460 149.870 132.660 150.170 ;
        RECT 141.640 149.870 144.530 150.295 ;
        RECT 26.640 148.410 29.040 148.710 ;
        RECT 26.340 148.110 29.040 148.410 ;
        RECT 34.230 148.575 34.680 149.300 ;
        RECT 44.195 149.025 47.405 149.445 ;
        RECT 43.605 148.855 47.405 149.025 ;
        RECT 43.605 148.575 46.795 148.855 ;
        RECT 34.230 148.255 46.795 148.575 ;
        RECT 34.230 148.125 46.195 148.255 ;
        RECT 25.740 147.510 29.640 148.110 ;
        RECT 43.030 147.755 46.195 148.125 ;
        RECT 42.460 147.645 46.195 147.755 ;
        RECT 15.085 147.080 17.495 147.500 ;
        RECT 14.685 146.695 17.495 147.080 ;
        RECT 14.685 146.265 17.085 146.695 ;
        RECT 14.295 145.890 17.085 146.265 ;
        RECT 25.440 146.310 29.940 147.510 ;
        RECT 42.460 147.105 45.605 147.645 ;
        RECT 41.905 147.025 45.605 147.105 ;
        RECT 41.905 146.445 45.030 147.025 ;
        RECT 25.440 146.010 26.340 146.310 ;
        RECT 14.295 145.445 16.685 145.890 ;
        RECT 25.440 145.710 26.040 146.010 ;
        RECT 13.915 145.080 16.685 145.445 ;
        RECT 25.740 145.410 26.040 145.710 ;
        RECT 27.240 145.410 28.140 146.310 ;
        RECT 29.040 146.010 29.940 146.310 ;
        RECT 29.340 145.710 29.940 146.010 ;
        RECT 41.360 146.395 45.030 146.445 ;
        RECT 41.360 145.775 44.460 146.395 ;
        RECT 40.830 145.755 44.460 145.775 ;
        RECT 29.340 145.410 29.640 145.710 ;
        RECT 25.740 145.110 26.340 145.410 ;
        RECT 26.940 145.110 28.440 145.410 ;
        RECT 29.040 145.110 29.640 145.410 ;
        RECT 13.915 144.615 16.295 145.080 ;
        RECT 25.740 144.810 27.540 145.110 ;
        RECT 27.840 144.810 29.340 145.110 ;
        RECT 40.830 145.105 43.905 145.755 ;
        RECT 40.830 145.095 43.360 145.105 ;
        RECT 13.545 144.265 16.295 144.615 ;
        RECT 26.340 144.510 27.240 144.810 ;
        RECT 28.140 144.510 29.340 144.810 ;
        RECT 13.545 143.785 15.915 144.265 ;
        RECT 26.640 143.910 28.740 144.510 ;
        RECT 40.310 144.445 43.360 145.095 ;
        RECT 40.310 144.410 42.830 144.445 ;
        RECT 13.185 143.445 15.915 143.785 ;
        RECT 24.840 143.610 25.740 143.910 ;
        RECT 26.640 143.610 26.940 143.910 ;
        RECT 27.240 143.610 27.540 143.910 ;
        RECT 27.840 143.610 28.140 143.910 ;
        RECT 28.440 143.610 28.740 143.910 ;
        RECT 29.640 143.610 30.540 143.910 ;
        RECT 39.800 143.775 42.830 144.410 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 112.855 149.445 116.685 149.645 ;
        RECT 113.475 149.025 116.685 149.445 ;
        RECT 130.560 149.270 132.060 149.870 ;
        RECT 142.090 149.500 144.530 149.870 ;
        RECT 113.475 148.855 117.275 149.025 ;
        RECT 129.960 148.970 131.160 149.270 ;
        RECT 131.460 148.970 132.660 149.270 ;
        RECT 142.090 149.085 144.960 149.500 ;
        RECT 114.085 148.395 117.275 148.855 ;
        RECT 128.460 148.670 130.560 148.970 ;
        RECT 132.060 148.670 134.460 148.970 ;
        RECT 114.085 148.255 117.850 148.395 ;
        RECT 114.685 147.755 117.850 148.255 ;
        RECT 128.160 148.370 129.960 148.670 ;
        RECT 132.660 148.370 134.460 148.670 ;
        RECT 128.160 148.070 129.360 148.370 ;
        RECT 133.260 148.070 134.460 148.370 ;
        RECT 142.530 148.695 144.960 149.085 ;
        RECT 142.530 148.295 145.385 148.695 ;
        RECT 128.160 147.770 129.060 148.070 ;
        RECT 133.560 147.770 134.460 148.070 ;
        RECT 142.960 147.890 145.385 148.295 ;
        RECT 114.685 147.645 118.420 147.755 ;
        RECT 115.275 147.105 118.420 147.645 ;
        RECT 128.460 147.470 128.760 147.770 ;
        RECT 130.260 147.470 130.560 147.770 ;
        RECT 130.860 147.470 131.160 147.770 ;
        RECT 131.460 147.470 131.760 147.770 ;
        RECT 132.060 147.470 132.360 147.770 ;
        RECT 133.860 147.470 134.160 147.770 ;
        RECT 142.960 147.500 145.795 147.890 ;
        RECT 115.275 147.025 118.975 147.105 ;
        RECT 115.850 146.445 118.975 147.025 ;
        RECT 130.260 146.870 132.360 147.470 ;
        RECT 143.385 147.080 145.795 147.500 ;
        RECT 129.960 146.570 130.860 146.870 ;
        RECT 131.760 146.570 132.960 146.870 ;
        RECT 143.385 146.695 146.195 147.080 ;
        RECT 115.850 146.395 119.520 146.445 ;
        RECT 116.420 145.775 119.520 146.395 ;
        RECT 129.360 146.270 131.160 146.570 ;
        RECT 131.460 146.270 132.960 146.570 ;
        RECT 129.360 145.970 129.960 146.270 ;
        RECT 130.560 145.970 132.060 146.270 ;
        RECT 132.660 145.970 133.260 146.270 ;
        RECT 116.420 145.755 120.050 145.775 ;
        RECT 116.975 145.105 120.050 145.755 ;
        RECT 129.360 145.670 129.660 145.970 ;
        RECT 117.520 145.095 120.050 145.105 ;
        RECT 129.060 145.370 129.660 145.670 ;
        RECT 117.520 144.445 120.570 145.095 ;
        RECT 118.050 144.410 120.570 144.445 ;
        RECT 129.060 145.070 129.960 145.370 ;
        RECT 130.860 145.070 131.760 145.970 ;
        RECT 132.960 145.670 133.260 145.970 ;
        RECT 143.795 146.265 146.195 146.695 ;
        RECT 143.795 145.890 146.585 146.265 ;
        RECT 132.960 145.370 133.560 145.670 ;
        RECT 132.660 145.070 133.560 145.370 ;
        RECT 144.195 145.445 146.585 145.890 ;
        RECT 144.195 145.080 146.965 145.445 ;
        RECT 39.800 143.715 42.310 143.775 ;
        RECT 13.185 142.950 15.545 143.445 ;
        RECT 24.540 143.010 26.040 143.610 ;
        RECT 29.340 143.010 30.840 143.610 ;
        RECT 39.305 143.095 42.310 143.715 ;
        RECT 39.305 143.010 41.800 143.095 ;
        RECT 12.835 142.615 15.545 142.950 ;
        RECT 24.840 142.710 26.640 143.010 ;
        RECT 28.740 142.710 30.540 143.010 ;
        RECT 12.835 142.110 15.185 142.615 ;
        RECT 25.740 142.410 26.940 142.710 ;
        RECT 28.440 142.410 29.640 142.710 ;
        RECT 38.820 142.410 41.800 143.010 ;
        RECT 26.340 142.110 27.540 142.410 ;
        RECT 27.840 142.110 29.040 142.410 ;
        RECT 38.820 142.295 41.305 142.410 ;
        RECT 12.500 141.785 15.185 142.110 ;
        RECT 12.500 141.270 14.835 141.785 ;
        RECT 26.940 141.510 28.440 142.110 ;
        RECT 38.350 141.715 41.305 142.295 ;
        RECT 38.350 141.575 40.820 141.715 ;
        RECT 12.170 140.950 14.835 141.270 ;
        RECT 26.340 141.210 27.540 141.510 ;
        RECT 27.840 141.210 29.040 141.510 ;
        RECT 12.170 140.420 14.500 140.950 ;
        RECT 24.840 140.910 26.940 141.210 ;
        RECT 28.440 140.910 30.840 141.210 ;
        RECT 11.855 140.110 14.500 140.420 ;
        RECT 24.540 140.610 26.340 140.910 ;
        RECT 29.040 140.610 30.840 140.910 ;
        RECT 37.890 141.010 40.820 141.575 ;
        RECT 37.890 140.845 40.350 141.010 ;
        RECT 24.540 140.310 25.740 140.610 ;
        RECT 29.640 140.310 30.840 140.610 ;
        RECT 11.855 139.570 14.170 140.110 ;
        RECT 24.540 140.010 25.440 140.310 ;
        RECT 29.940 140.010 30.840 140.310 ;
        RECT 37.440 140.295 40.350 140.845 ;
        RECT 37.440 140.105 39.890 140.295 ;
        RECT 24.840 139.710 25.140 140.010 ;
        RECT 26.640 139.710 26.940 140.010 ;
        RECT 27.240 139.710 27.540 140.010 ;
        RECT 27.840 139.710 28.140 140.010 ;
        RECT 28.440 139.710 28.740 140.010 ;
        RECT 30.240 139.710 30.540 140.010 ;
        RECT 11.545 139.270 14.170 139.570 ;
        RECT 11.545 138.715 13.855 139.270 ;
        RECT 26.640 139.110 28.740 139.710 ;
        RECT 37.005 139.575 39.890 140.105 ;
        RECT 37.005 139.365 39.440 139.575 ;
        RECT 26.340 138.810 27.240 139.110 ;
        RECT 28.140 138.810 29.340 139.110 ;
        RECT 11.250 138.420 13.855 138.715 ;
        RECT 25.740 138.510 27.540 138.810 ;
        RECT 27.840 138.510 29.340 138.810 ;
        RECT 36.585 138.845 39.440 139.365 ;
        RECT 36.585 138.610 39.005 138.845 ;
        RECT 11.250 137.855 13.545 138.420 ;
        RECT 25.740 138.210 26.340 138.510 ;
        RECT 26.940 138.210 28.440 138.510 ;
        RECT 29.040 138.210 29.640 138.510 ;
        RECT 25.740 137.910 26.040 138.210 ;
        RECT 10.965 137.570 13.545 137.855 ;
        RECT 25.440 137.610 26.040 137.910 ;
        RECT 10.965 136.995 13.250 137.570 ;
        RECT 10.690 136.715 13.250 136.995 ;
        RECT 25.440 137.310 26.340 137.610 ;
        RECT 27.240 137.310 28.140 138.210 ;
        RECT 29.340 137.910 29.640 138.210 ;
        RECT 36.180 138.105 39.005 138.610 ;
        RECT 29.340 137.610 29.940 137.910 ;
        RECT 36.180 137.855 38.585 138.105 ;
        RECT 29.040 137.310 29.940 137.610 ;
        RECT 10.690 136.130 12.965 136.715 ;
        RECT 10.430 135.855 12.965 136.130 ;
        RECT 25.440 136.110 29.940 137.310 ;
        RECT 35.785 137.365 38.585 137.855 ;
        RECT 35.785 137.090 38.180 137.365 ;
        RECT 35.400 136.610 38.180 137.090 ;
        RECT 35.400 136.315 37.785 136.610 ;
        RECT 10.430 135.260 12.690 135.855 ;
        RECT 10.175 134.995 12.690 135.260 ;
        RECT 10.175 134.390 12.430 134.995 ;
        RECT 9.935 134.130 12.430 134.390 ;
        RECT 24.160 134.520 24.720 135.910 ;
        RECT 25.740 135.510 29.640 136.110 ;
        RECT 35.035 135.855 37.785 136.315 ;
        RECT 35.035 135.540 37.400 135.855 ;
        RECT 26.340 135.210 29.040 135.510 ;
        RECT 26.640 134.910 29.040 135.210 ;
        RECT 34.680 135.090 37.400 135.540 ;
        RECT 34.680 134.755 37.035 135.090 ;
        RECT 9.935 133.515 12.175 134.130 ;
        RECT 24.160 134.090 24.610 134.520 ;
        RECT 34.340 134.315 37.035 134.755 ;
        RECT 34.340 134.090 36.680 134.315 ;
        RECT 24.160 133.640 36.680 134.090 ;
        RECT 9.705 133.260 12.175 133.515 ;
        RECT 34.010 133.540 36.680 133.640 ;
        RECT 60.370 134.000 99.370 144.400 ;
        RECT 118.050 143.775 121.080 144.410 ;
        RECT 129.060 143.870 133.560 145.070 ;
        RECT 144.585 144.615 146.965 145.080 ;
        RECT 144.585 144.265 147.335 144.615 ;
        RECT 118.570 143.715 121.080 143.775 ;
        RECT 118.570 143.095 121.575 143.715 ;
        RECT 119.080 143.010 121.575 143.095 ;
        RECT 119.080 142.410 122.060 143.010 ;
        RECT 119.575 142.295 122.060 142.410 ;
        RECT 119.575 141.850 122.530 142.295 ;
        RECT 127.780 142.280 128.340 143.670 ;
        RECT 129.360 143.270 133.260 143.870 ;
        RECT 144.965 143.785 147.335 144.265 ;
        RECT 144.965 143.445 147.695 143.785 ;
        RECT 129.960 142.970 132.660 143.270 ;
        RECT 130.260 142.670 132.660 142.970 ;
        RECT 145.335 142.950 147.695 143.445 ;
        RECT 145.335 142.615 148.045 142.950 ;
        RECT 127.780 141.850 128.230 142.280 ;
        RECT 119.575 141.715 128.230 141.850 ;
        RECT 145.695 142.110 148.045 142.615 ;
        RECT 145.695 141.785 148.380 142.110 ;
        RECT 120.060 141.400 128.230 141.715 ;
        RECT 120.060 141.010 122.990 141.400 ;
        RECT 146.045 141.290 148.380 141.785 ;
        RECT 120.530 140.845 122.990 141.010 ;
        RECT 139.550 141.270 148.380 141.290 ;
        RECT 120.530 140.295 123.440 140.845 ;
        RECT 139.550 140.840 148.710 141.270 ;
        RECT 120.990 140.105 123.440 140.295 ;
        RECT 120.990 139.575 123.875 140.105 ;
        RECT 135.120 140.060 137.520 140.360 ;
        RECT 135.120 139.760 137.820 140.060 ;
        RECT 121.440 139.365 123.875 139.575 ;
        RECT 121.440 138.845 124.295 139.365 ;
        RECT 134.520 139.160 138.420 139.760 ;
        RECT 139.550 139.290 140.000 140.840 ;
        RECT 146.380 140.420 148.710 140.840 ;
        RECT 146.380 140.110 149.025 140.420 ;
        RECT 146.710 139.570 149.025 140.110 ;
        RECT 146.710 139.270 149.335 139.570 ;
        RECT 121.875 138.610 124.295 138.845 ;
        RECT 121.875 138.105 124.700 138.610 ;
        RECT 122.295 137.855 124.700 138.105 ;
        RECT 134.220 137.960 138.720 139.160 ;
        RECT 147.025 138.715 149.335 139.270 ;
        RECT 147.025 138.420 149.630 138.715 ;
        RECT 122.295 137.365 125.095 137.855 ;
        RECT 122.700 137.090 125.095 137.365 ;
        RECT 134.220 137.660 135.120 137.960 ;
        RECT 134.220 137.360 134.820 137.660 ;
        RECT 122.700 136.610 125.480 137.090 ;
        RECT 134.520 137.060 134.820 137.360 ;
        RECT 136.020 137.060 136.920 137.960 ;
        RECT 137.820 137.660 138.720 137.960 ;
        RECT 138.120 137.360 138.720 137.660 ;
        RECT 147.335 137.855 149.630 138.420 ;
        RECT 147.335 137.570 149.915 137.855 ;
        RECT 138.120 137.060 138.420 137.360 ;
        RECT 134.520 136.760 135.120 137.060 ;
        RECT 135.720 136.760 137.220 137.060 ;
        RECT 137.820 136.760 138.420 137.060 ;
        RECT 123.095 136.315 125.480 136.610 ;
        RECT 134.820 136.460 136.320 136.760 ;
        RECT 136.620 136.460 138.420 136.760 ;
        RECT 147.630 136.995 149.915 137.570 ;
        RECT 147.630 136.715 150.190 136.995 ;
        RECT 123.095 135.855 125.845 136.315 ;
        RECT 134.820 136.160 136.020 136.460 ;
        RECT 136.920 136.160 137.820 136.460 ;
        RECT 123.480 135.540 125.845 135.855 ;
        RECT 135.420 135.560 137.520 136.160 ;
        RECT 147.915 136.130 150.190 136.715 ;
        RECT 147.915 135.855 150.450 136.130 ;
        RECT 123.480 135.090 126.200 135.540 ;
        RECT 133.620 135.260 134.520 135.560 ;
        RECT 135.420 135.260 135.720 135.560 ;
        RECT 136.020 135.260 136.320 135.560 ;
        RECT 136.620 135.260 136.920 135.560 ;
        RECT 137.220 135.260 137.520 135.560 ;
        RECT 138.420 135.260 139.320 135.560 ;
        RECT 148.190 135.260 150.450 135.855 ;
        RECT 123.845 134.755 126.200 135.090 ;
        RECT 123.845 134.315 126.540 134.755 ;
        RECT 133.320 134.660 134.820 135.260 ;
        RECT 138.120 134.660 139.620 135.260 ;
        RECT 148.190 134.995 150.705 135.260 ;
        RECT 133.620 134.360 135.420 134.660 ;
        RECT 137.520 134.360 139.320 134.660 ;
        RECT 148.450 134.390 150.705 134.995 ;
        RECT 9.705 132.635 11.935 133.260 ;
        RECT 34.010 133.170 36.340 133.540 ;
        RECT 9.485 132.505 11.935 132.635 ;
        RECT 33.695 132.755 36.340 133.170 ;
        RECT 22.900 132.505 23.350 132.550 ;
        RECT 9.485 132.055 23.350 132.505 ;
        RECT 33.695 132.365 36.010 132.755 ;
        RECT 9.485 131.755 11.705 132.055 ;
        RECT 9.275 131.515 11.705 131.755 ;
        RECT 9.275 130.870 11.485 131.515 ;
        RECT 18.470 131.320 20.870 131.620 ;
        RECT 18.470 131.020 21.170 131.320 ;
        RECT 9.080 130.635 11.485 130.870 ;
        RECT 9.080 129.985 11.275 130.635 ;
        RECT 17.870 130.420 21.770 131.020 ;
        RECT 22.900 130.550 23.350 132.055 ;
        RECT 33.400 131.965 36.010 132.365 ;
        RECT 33.400 131.560 35.695 131.965 ;
        RECT 33.110 131.170 35.695 131.560 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 33.110 130.750 35.400 131.170 ;
        RECT 8.895 129.755 11.275 129.985 ;
        RECT 8.895 129.100 11.080 129.755 ;
        RECT 8.720 128.870 11.080 129.100 ;
        RECT 17.570 129.220 22.070 130.420 ;
        RECT 32.840 130.365 35.400 130.750 ;
        RECT 32.840 129.935 35.110 130.365 ;
        RECT 17.570 128.920 18.470 129.220 ;
        RECT 8.720 128.210 10.895 128.870 ;
        RECT 17.570 128.620 18.170 128.920 ;
        RECT 8.555 127.985 10.895 128.210 ;
        RECT 17.870 128.320 18.170 128.620 ;
        RECT 19.370 128.320 20.270 129.220 ;
        RECT 21.170 128.920 22.070 129.220 ;
        RECT 32.585 129.560 35.110 129.935 ;
        RECT 32.585 129.115 34.840 129.560 ;
        RECT 21.470 128.620 22.070 128.920 ;
        RECT 32.340 128.750 34.840 129.115 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 21.470 128.320 21.770 128.620 ;
        RECT 17.870 128.020 18.470 128.320 ;
        RECT 19.070 128.020 20.570 128.320 ;
        RECT 21.170 128.020 21.770 128.320 ;
        RECT 32.340 128.290 34.585 128.750 ;
        RECT 8.555 127.315 10.720 127.985 ;
        RECT 18.170 127.720 19.670 128.020 ;
        RECT 19.970 127.720 21.770 128.020 ;
        RECT 32.110 127.935 34.585 128.290 ;
        RECT 18.170 127.420 19.370 127.720 ;
        RECT 20.270 127.420 21.170 127.720 ;
        RECT 32.110 127.460 34.340 127.935 ;
        RECT 8.400 127.100 10.720 127.315 ;
        RECT 8.400 126.425 10.555 127.100 ;
        RECT 18.770 126.820 20.870 127.420 ;
        RECT 31.900 127.115 34.340 127.460 ;
        RECT 16.970 126.520 17.870 126.820 ;
        RECT 18.770 126.520 19.070 126.820 ;
        RECT 19.370 126.520 19.670 126.820 ;
        RECT 19.970 126.520 20.270 126.820 ;
        RECT 20.570 126.520 20.870 126.820 ;
        RECT 21.770 126.520 22.670 126.820 ;
        RECT 31.900 126.630 34.110 127.115 ;
        RECT 8.260 126.210 10.555 126.425 ;
        RECT 8.260 125.530 10.400 126.210 ;
        RECT 16.670 125.920 18.170 126.520 ;
        RECT 21.470 125.920 22.970 126.520 ;
        RECT 31.700 126.290 34.110 126.630 ;
        RECT 16.970 125.620 18.770 125.920 ;
        RECT 20.870 125.620 22.670 125.920 ;
        RECT 31.700 125.795 33.900 126.290 ;
        RECT 8.130 125.315 10.400 125.530 ;
        RECT 17.870 125.320 19.070 125.620 ;
        RECT 20.570 125.320 21.770 125.620 ;
        RECT 31.515 125.460 33.900 125.795 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 124.200 133.965 126.540 134.315 ;
        RECT 134.520 134.060 135.720 134.360 ;
        RECT 137.220 134.060 138.420 134.360 ;
        RECT 148.450 134.130 150.945 134.390 ;
        RECT 124.200 133.540 126.870 133.965 ;
        RECT 135.120 133.760 136.320 134.060 ;
        RECT 136.620 133.760 137.820 134.060 ;
        RECT 124.540 133.170 126.870 133.540 ;
        RECT 124.540 132.755 127.185 133.170 ;
        RECT 135.720 133.160 137.220 133.760 ;
        RECT 148.705 133.515 150.945 134.130 ;
        RECT 148.705 133.260 151.175 133.515 ;
        RECT 135.120 132.860 136.320 133.160 ;
        RECT 136.620 132.860 137.820 133.160 ;
        RECT 124.870 132.365 127.185 132.755 ;
        RECT 133.320 132.560 135.720 132.860 ;
        RECT 137.220 132.560 139.320 132.860 ;
        RECT 148.945 132.635 151.175 133.260 ;
        RECT 124.870 131.965 127.480 132.365 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 125.185 131.560 127.480 131.965 ;
        RECT 133.320 132.260 135.120 132.560 ;
        RECT 137.820 132.260 139.620 132.560 ;
        RECT 148.945 132.390 151.395 132.635 ;
        RECT 133.320 131.960 134.520 132.260 ;
        RECT 138.420 131.960 139.620 132.260 ;
        RECT 133.320 131.660 134.220 131.960 ;
        RECT 138.720 131.660 139.620 131.960 ;
        RECT 149.175 131.755 151.395 132.390 ;
        RECT 125.185 131.170 127.770 131.560 ;
        RECT 133.620 131.360 133.920 131.660 ;
        RECT 135.420 131.360 135.720 131.660 ;
        RECT 136.020 131.360 136.320 131.660 ;
        RECT 136.620 131.360 136.920 131.660 ;
        RECT 137.220 131.360 137.520 131.660 ;
        RECT 139.020 131.360 139.320 131.660 ;
        RECT 149.175 131.515 151.605 131.755 ;
        RECT 125.480 130.750 127.770 131.170 ;
        RECT 135.420 130.760 137.520 131.360 ;
        RECT 149.395 130.870 151.605 131.515 ;
        RECT 125.480 130.365 128.040 130.750 ;
        RECT 125.770 129.935 128.040 130.365 ;
        RECT 134.820 130.460 136.020 130.760 ;
        RECT 136.920 130.460 137.820 130.760 ;
        RECT 149.395 130.635 151.800 130.870 ;
        RECT 134.820 130.160 136.320 130.460 ;
        RECT 136.620 130.160 138.420 130.460 ;
        RECT 125.770 129.560 128.295 129.935 ;
        RECT 134.520 129.860 135.120 130.160 ;
        RECT 135.720 129.860 137.220 130.160 ;
        RECT 137.820 129.860 138.420 130.160 ;
        RECT 134.520 129.560 134.820 129.860 ;
        RECT 126.040 129.115 128.295 129.560 ;
        RECT 134.220 129.260 134.820 129.560 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 126.040 128.750 128.540 129.115 ;
        RECT 126.295 128.290 128.540 128.750 ;
        RECT 134.220 128.960 135.120 129.260 ;
        RECT 136.020 128.960 136.920 129.860 ;
        RECT 138.120 129.560 138.420 129.860 ;
        RECT 149.605 129.985 151.800 130.635 ;
        RECT 149.605 129.755 151.985 129.985 ;
        RECT 138.120 129.260 138.720 129.560 ;
        RECT 137.820 128.960 138.720 129.260 ;
        RECT 126.295 127.935 128.770 128.290 ;
        RECT 126.540 127.460 128.770 127.935 ;
        RECT 134.220 127.760 138.720 128.960 ;
        RECT 149.800 129.100 151.985 129.755 ;
        RECT 149.800 128.870 152.160 129.100 ;
        RECT 149.985 128.210 152.160 128.870 ;
        RECT 149.985 127.985 152.325 128.210 ;
        RECT 126.540 127.115 128.980 127.460 ;
        RECT 134.520 127.160 138.420 127.760 ;
        RECT 126.770 126.630 128.980 127.115 ;
        RECT 135.120 126.860 137.820 127.160 ;
        RECT 126.770 126.290 129.180 126.630 ;
        RECT 135.120 126.560 137.520 126.860 ;
        RECT 8.130 124.630 10.260 125.315 ;
        RECT 18.470 125.020 19.670 125.320 ;
        RECT 19.970 125.020 21.170 125.320 ;
        RECT 8.010 124.425 10.260 124.630 ;
        RECT 8.010 123.735 10.130 124.425 ;
        RECT 19.070 124.420 20.570 125.020 ;
        RECT 31.515 124.955 33.700 125.460 ;
        RECT 31.345 124.630 33.700 124.955 ;
        RECT 18.470 124.120 19.670 124.420 ;
        RECT 19.970 124.120 21.170 124.420 ;
        RECT 7.900 123.530 10.130 123.735 ;
        RECT 16.670 123.820 19.070 124.120 ;
        RECT 20.570 123.820 22.670 124.120 ;
        RECT 31.345 124.115 33.515 124.630 ;
        RECT 7.900 122.835 10.010 123.530 ;
        RECT 16.670 123.520 18.470 123.820 ;
        RECT 21.170 123.520 22.970 123.820 ;
        RECT 16.670 123.220 17.870 123.520 ;
        RECT 21.770 123.220 22.970 123.520 ;
        RECT 31.185 123.795 33.515 124.115 ;
        RECT 31.185 123.275 33.345 123.795 ;
        RECT 16.670 122.920 17.570 123.220 ;
        RECT 22.070 122.920 22.970 123.220 ;
        RECT 31.045 122.955 33.345 123.275 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
        RECT 126.980 125.795 129.180 126.290 ;
        RECT 139.440 126.170 140.000 127.560 ;
        RECT 150.160 127.315 152.325 127.985 ;
        RECT 150.160 127.100 152.480 127.315 ;
        RECT 150.325 126.425 152.480 127.100 ;
        RECT 150.325 126.210 152.620 126.425 ;
        RECT 126.980 125.740 129.365 125.795 ;
        RECT 139.550 125.740 140.000 126.170 ;
        RECT 126.980 125.460 140.000 125.740 ;
        RECT 127.180 125.290 140.000 125.460 ;
        RECT 150.480 125.530 152.620 126.210 ;
        RECT 150.480 125.315 152.750 125.530 ;
        RECT 127.180 124.955 129.365 125.290 ;
        RECT 127.180 124.630 129.535 124.955 ;
        RECT 127.365 124.115 129.535 124.630 ;
        RECT 150.620 124.630 152.750 125.315 ;
        RECT 150.620 124.425 152.870 124.630 ;
        RECT 127.365 123.795 129.695 124.115 ;
        RECT 7.805 122.630 10.010 122.835 ;
        RECT 7.805 121.935 9.900 122.630 ;
        RECT 16.970 122.620 17.270 122.920 ;
        RECT 18.770 122.620 19.070 122.920 ;
        RECT 19.370 122.620 19.670 122.920 ;
        RECT 19.970 122.620 20.270 122.920 ;
        RECT 20.570 122.620 20.870 122.920 ;
        RECT 22.370 122.620 22.670 122.920 ;
        RECT 18.770 122.020 20.870 122.620 ;
        RECT 31.045 122.425 33.185 122.955 ;
        RECT 30.920 122.115 33.185 122.425 ;
        RECT 7.720 121.735 9.900 121.935 ;
        RECT 7.720 121.030 9.805 121.735 ;
        RECT 18.170 121.720 19.370 122.020 ;
        RECT 20.270 121.720 21.170 122.020 ;
        RECT 18.170 121.420 19.670 121.720 ;
        RECT 19.970 121.420 21.770 121.720 ;
        RECT 30.920 121.580 33.045 122.115 ;
        RECT 7.645 120.835 9.805 121.030 ;
        RECT 17.870 121.120 18.470 121.420 ;
        RECT 19.070 121.120 20.570 121.420 ;
        RECT 21.170 121.120 21.770 121.420 ;
        RECT 7.645 120.130 9.720 120.835 ;
        RECT 17.870 120.820 18.170 121.120 ;
        RECT 7.585 119.935 9.720 120.130 ;
        RECT 17.570 120.520 18.170 120.820 ;
        RECT 17.570 120.220 18.470 120.520 ;
        RECT 19.370 120.220 20.270 121.120 ;
        RECT 21.470 120.820 21.770 121.120 ;
        RECT 30.810 121.275 33.045 121.580 ;
        RECT 21.470 120.520 22.070 120.820 ;
        RECT 30.810 120.730 32.920 121.275 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 127.535 123.275 129.695 123.795 ;
        RECT 150.750 123.735 152.870 124.425 ;
        RECT 150.750 123.610 152.980 123.735 ;
        RECT 127.535 122.955 129.835 123.275 ;
        RECT 127.695 122.425 129.835 122.955 ;
        RECT 138.210 123.160 152.980 123.610 ;
        RECT 127.695 122.115 129.960 122.425 ;
        RECT 127.835 121.580 129.960 122.115 ;
        RECT 138.210 121.610 138.660 123.160 ;
        RECT 150.870 122.835 152.980 123.160 ;
        RECT 140.690 122.380 143.090 122.680 ;
        RECT 150.870 122.630 153.075 122.835 ;
        RECT 140.390 122.080 143.090 122.380 ;
        RECT 127.835 121.275 130.070 121.580 ;
        RECT 139.790 121.480 143.690 122.080 ;
        RECT 150.980 121.935 153.075 122.630 ;
        RECT 150.980 121.735 153.160 121.935 ;
        RECT 21.170 120.220 22.070 120.520 ;
        RECT 7.585 119.225 9.645 119.935 ;
        RECT 7.535 119.030 9.645 119.225 ;
        RECT 7.535 118.320 9.585 119.030 ;
        RECT 17.570 119.020 22.070 120.220 ;
        RECT 30.710 120.425 32.920 120.730 ;
        RECT 30.710 119.880 32.810 120.425 ;
        RECT 30.630 119.580 32.810 119.880 ;
        RECT 30.630 119.025 32.710 119.580 ;
        RECT 17.870 118.420 21.770 119.020 ;
        RECT 7.495 118.130 9.585 118.320 ;
        RECT 7.495 117.415 9.535 118.130 ;
        RECT 18.470 118.120 21.170 118.420 ;
        RECT 18.470 117.820 20.870 118.120 ;
        RECT 22.790 117.430 23.350 118.820 ;
        RECT 30.560 118.730 32.710 119.025 ;
        RECT 30.560 118.170 32.630 118.730 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 127.960 120.730 130.070 121.275 ;
        RECT 127.960 120.425 130.170 120.730 ;
        RECT 128.070 119.880 130.170 120.425 ;
        RECT 139.490 120.280 143.990 121.480 ;
        RECT 151.075 121.030 153.160 121.735 ;
        RECT 151.075 120.835 153.235 121.030 ;
        RECT 139.490 119.980 140.390 120.280 ;
        RECT 128.070 119.580 130.250 119.880 ;
        RECT 139.490 119.680 140.090 119.980 ;
        RECT 128.170 119.025 130.250 119.580 ;
        RECT 139.790 119.380 140.090 119.680 ;
        RECT 141.290 119.380 142.190 120.280 ;
        RECT 143.090 119.980 143.990 120.280 ;
        RECT 143.390 119.680 143.990 119.980 ;
        RECT 151.160 120.130 153.235 120.835 ;
        RECT 151.160 119.935 153.295 120.130 ;
        RECT 143.390 119.380 143.690 119.680 ;
        RECT 139.790 119.080 140.390 119.380 ;
        RECT 140.990 119.080 142.490 119.380 ;
        RECT 143.090 119.080 143.690 119.380 ;
        RECT 151.235 119.225 153.295 119.935 ;
        RECT 128.170 118.730 130.320 119.025 ;
        RECT 139.790 118.780 141.590 119.080 ;
        RECT 141.890 118.780 143.390 119.080 ;
        RECT 151.235 119.030 153.345 119.225 ;
        RECT 7.465 117.225 9.535 117.415 ;
        RECT 7.465 116.510 9.495 117.225 ;
        RECT 22.900 117.045 23.350 117.430 ;
        RECT 30.510 117.880 32.630 118.170 ;
        RECT 30.510 117.320 32.560 117.880 ;
        RECT 30.470 117.045 32.560 117.320 ;
        RECT 22.900 117.025 32.560 117.045 ;
        RECT 22.900 116.595 32.510 117.025 ;
        RECT 22.900 116.550 23.350 116.595 ;
        RECT 7.450 116.320 9.495 116.510 ;
        RECT 7.450 115.610 9.465 116.320 ;
        RECT 30.450 116.170 32.510 116.595 ;
        RECT 30.450 115.610 32.470 116.170 ;
        RECT 7.440 115.415 9.465 115.610 ;
        RECT 7.440 114.670 9.450 115.415 ;
        RECT 30.440 115.320 32.470 115.610 ;
        RECT 7.440 114.220 19.340 114.670 ;
        RECT 7.440 113.805 9.450 114.220 ;
        RECT 7.440 113.615 9.465 113.805 ;
        RECT 7.450 112.900 9.465 113.615 ;
        RECT 7.450 112.710 9.495 112.900 ;
        RECT 7.465 111.995 9.495 112.710 ;
        RECT 18.890 112.670 19.340 114.220 ;
        RECT 30.440 113.900 32.450 115.320 ;
        RECT 21.370 113.440 23.770 113.740 ;
        RECT 30.440 113.615 32.470 113.900 ;
        RECT 21.070 113.140 23.770 113.440 ;
        RECT 20.470 112.540 24.370 113.140 ;
        RECT 30.450 113.050 32.470 113.615 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 128.250 118.170 130.320 118.730 ;
        RECT 140.390 118.480 141.290 118.780 ;
        RECT 142.190 118.480 143.390 118.780 ;
        RECT 128.250 117.880 130.370 118.170 ;
        RECT 140.690 117.880 142.790 118.480 ;
        RECT 151.295 118.320 153.345 119.030 ;
        RECT 151.295 118.130 153.385 118.320 ;
        RECT 128.320 117.320 130.370 117.880 ;
        RECT 138.890 117.580 139.790 117.880 ;
        RECT 140.690 117.580 140.990 117.880 ;
        RECT 141.290 117.580 141.590 117.880 ;
        RECT 141.890 117.580 142.190 117.880 ;
        RECT 142.490 117.580 142.790 117.880 ;
        RECT 143.690 117.580 144.590 117.880 ;
        RECT 128.320 117.025 130.410 117.320 ;
        RECT 128.370 116.465 130.410 117.025 ;
        RECT 138.590 116.980 140.090 117.580 ;
        RECT 143.390 116.980 144.890 117.580 ;
        RECT 151.345 117.415 153.385 118.130 ;
        RECT 151.345 117.225 153.415 117.415 ;
        RECT 138.890 116.680 140.690 116.980 ;
        RECT 142.790 116.680 144.590 116.980 ;
        RECT 128.370 116.170 130.430 116.465 ;
        RECT 139.790 116.380 140.990 116.680 ;
        RECT 142.490 116.380 143.690 116.680 ;
        RECT 151.385 116.510 153.415 117.225 ;
        RECT 128.410 115.610 130.430 116.170 ;
        RECT 140.390 116.080 141.590 116.380 ;
        RECT 141.890 116.080 143.090 116.380 ;
        RECT 151.385 116.320 153.430 116.510 ;
        RECT 128.410 115.320 130.440 115.610 ;
        RECT 140.990 115.480 142.490 116.080 ;
        RECT 151.415 115.610 153.430 116.320 ;
        RECT 128.430 113.900 130.440 115.320 ;
        RECT 140.390 115.180 141.590 115.480 ;
        RECT 141.890 115.180 143.090 115.480 ;
        RECT 151.415 115.415 153.440 115.610 ;
        RECT 138.890 114.880 140.990 115.180 ;
        RECT 142.490 114.880 144.890 115.180 ;
        RECT 138.590 114.580 140.390 114.880 ;
        RECT 143.090 114.580 144.890 114.880 ;
        RECT 138.590 114.280 139.790 114.580 ;
        RECT 143.690 114.280 144.890 114.580 ;
        RECT 138.590 113.980 139.490 114.280 ;
        RECT 143.990 113.980 144.890 114.280 ;
        RECT 128.410 113.610 130.440 113.900 ;
        RECT 138.890 113.680 139.190 113.980 ;
        RECT 140.690 113.680 140.990 113.980 ;
        RECT 141.290 113.680 141.590 113.980 ;
        RECT 141.890 113.680 142.190 113.980 ;
        RECT 142.490 113.680 142.790 113.980 ;
        RECT 144.290 113.680 144.590 113.980 ;
        RECT 151.430 113.805 153.440 115.415 ;
        RECT 30.450 112.755 32.510 113.050 ;
        RECT 7.465 111.805 9.535 111.995 ;
        RECT 7.495 111.090 9.535 111.805 ;
        RECT 20.170 111.340 24.670 112.540 ;
        RECT 30.470 112.195 32.510 112.755 ;
        RECT 30.470 111.900 32.560 112.195 ;
        RECT 7.495 110.900 9.585 111.090 ;
        RECT 7.535 110.190 9.585 110.900 ;
        RECT 20.170 111.040 21.070 111.340 ;
        RECT 20.170 110.740 20.770 111.040 ;
        RECT 20.470 110.440 20.770 110.740 ;
        RECT 21.970 110.440 22.870 111.340 ;
        RECT 23.770 111.040 24.670 111.340 ;
        RECT 30.510 111.340 32.560 111.900 ;
        RECT 30.510 111.050 32.630 111.340 ;
        RECT 24.070 110.740 24.670 111.040 ;
        RECT 24.070 110.440 24.370 110.740 ;
        RECT 7.535 109.995 9.645 110.190 ;
        RECT 7.585 109.285 9.645 109.995 ;
        RECT 20.470 110.140 21.070 110.440 ;
        RECT 21.670 110.140 23.170 110.440 ;
        RECT 23.770 110.140 24.370 110.440 ;
        RECT 30.560 110.490 32.630 111.050 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 128.410 113.050 130.430 113.610 ;
        RECT 140.690 113.080 142.790 113.680 ;
        RECT 151.415 113.610 153.440 113.805 ;
        RECT 128.370 112.755 130.430 113.050 ;
        RECT 140.390 112.780 141.290 113.080 ;
        RECT 142.190 112.780 143.390 113.080 ;
        RECT 151.415 112.900 153.430 113.610 ;
        RECT 128.370 112.195 130.410 112.755 ;
        RECT 128.320 111.900 130.410 112.195 ;
        RECT 139.790 112.480 141.590 112.780 ;
        RECT 141.890 112.480 143.390 112.780 ;
        RECT 151.385 112.710 153.430 112.900 ;
        RECT 139.790 112.180 140.390 112.480 ;
        RECT 140.990 112.180 142.490 112.480 ;
        RECT 143.090 112.180 143.690 112.480 ;
        RECT 128.320 111.340 130.370 111.900 ;
        RECT 139.790 111.880 140.090 112.180 ;
        RECT 128.250 111.050 130.370 111.340 ;
        RECT 139.490 111.580 140.090 111.880 ;
        RECT 139.490 111.280 140.390 111.580 ;
        RECT 141.290 111.280 142.190 112.180 ;
        RECT 143.390 111.880 143.690 112.180 ;
        RECT 151.385 111.995 153.415 112.710 ;
        RECT 143.390 111.580 143.990 111.880 ;
        RECT 143.090 111.280 143.990 111.580 ;
        RECT 30.560 110.195 32.710 110.490 ;
        RECT 20.470 109.840 22.270 110.140 ;
        RECT 22.570 109.840 24.070 110.140 ;
        RECT 21.070 109.540 21.970 109.840 ;
        RECT 22.870 109.540 24.070 109.840 ;
        RECT 30.630 109.640 32.710 110.195 ;
        RECT 7.585 109.090 9.720 109.285 ;
        RECT 7.645 108.385 9.720 109.090 ;
        RECT 21.370 108.940 23.470 109.540 ;
        RECT 30.630 109.340 32.810 109.640 ;
        RECT 19.570 108.640 20.470 108.940 ;
        RECT 21.370 108.640 21.670 108.940 ;
        RECT 21.970 108.640 22.270 108.940 ;
        RECT 22.570 108.640 22.870 108.940 ;
        RECT 23.170 108.640 23.470 108.940 ;
        RECT 24.370 108.640 25.270 108.940 ;
        RECT 30.710 108.795 32.810 109.340 ;
        RECT 7.645 108.190 9.805 108.385 ;
        RECT 7.720 107.485 9.805 108.190 ;
        RECT 19.270 108.040 20.770 108.640 ;
        RECT 24.070 108.040 25.570 108.640 ;
        RECT 30.710 108.490 32.920 108.795 ;
        RECT 19.570 107.740 21.370 108.040 ;
        RECT 23.470 107.740 25.270 108.040 ;
        RECT 30.810 107.945 32.920 108.490 ;
        RECT 7.720 107.285 9.900 107.485 ;
        RECT 20.470 107.440 21.670 107.740 ;
        RECT 23.170 107.440 24.370 107.740 ;
        RECT 30.810 107.640 33.045 107.945 ;
        RECT 7.805 106.590 9.900 107.285 ;
        RECT 21.070 107.140 22.270 107.440 ;
        RECT 22.570 107.140 23.770 107.440 ;
        RECT 7.805 106.385 10.010 106.590 ;
        RECT 21.670 106.540 23.170 107.140 ;
        RECT 30.920 107.105 33.045 107.640 ;
        RECT 30.920 106.795 33.185 107.105 ;
        RECT 7.900 105.690 10.010 106.385 ;
        RECT 21.070 106.240 22.270 106.540 ;
        RECT 22.570 106.240 23.770 106.540 ;
        RECT 31.045 106.265 33.185 106.795 ;
        RECT 19.570 105.940 21.670 106.240 ;
        RECT 23.170 105.940 25.570 106.240 ;
        RECT 31.045 105.945 33.345 106.265 ;
        RECT 7.900 105.485 10.130 105.690 ;
        RECT 8.010 104.795 10.130 105.485 ;
        RECT 19.270 105.640 21.070 105.940 ;
        RECT 23.770 105.640 25.570 105.940 ;
        RECT 19.270 105.340 20.470 105.640 ;
        RECT 24.370 105.340 25.570 105.640 ;
        RECT 19.270 105.040 20.170 105.340 ;
        RECT 24.670 105.040 25.570 105.340 ;
        RECT 31.185 105.425 33.345 105.945 ;
        RECT 31.185 105.105 33.515 105.425 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
        RECT 128.250 110.490 130.320 111.050 ;
        RECT 128.170 110.195 130.320 110.490 ;
        RECT 128.170 109.640 130.250 110.195 ;
        RECT 139.490 110.080 143.990 111.280 ;
        RECT 151.345 111.805 153.415 111.995 ;
        RECT 151.345 111.090 153.385 111.805 ;
        RECT 151.295 110.900 153.385 111.090 ;
        RECT 151.295 110.190 153.345 110.900 ;
        RECT 128.070 109.340 130.250 109.640 ;
        RECT 128.070 108.795 130.170 109.340 ;
        RECT 127.960 108.490 130.170 108.795 ;
        RECT 138.210 108.490 138.770 109.880 ;
        RECT 139.790 109.480 143.690 110.080 ;
        RECT 151.235 109.995 153.345 110.190 ;
        RECT 140.390 109.180 143.090 109.480 ;
        RECT 151.235 109.285 153.295 109.995 ;
        RECT 140.690 108.880 143.090 109.180 ;
        RECT 151.160 109.090 153.295 109.285 ;
        RECT 127.960 108.060 130.070 108.490 ;
        RECT 138.210 108.060 138.660 108.490 ;
        RECT 151.160 108.385 153.235 109.090 ;
        RECT 127.960 107.945 138.660 108.060 ;
        RECT 127.835 107.610 138.660 107.945 ;
        RECT 151.075 108.190 153.235 108.385 ;
        RECT 127.835 107.105 129.960 107.610 ;
        RECT 151.075 107.485 153.160 108.190 ;
        RECT 127.695 106.795 129.960 107.105 ;
        RECT 150.980 107.285 153.160 107.485 ;
        RECT 127.695 106.265 129.835 106.795 ;
        RECT 150.980 106.590 153.075 107.285 ;
        RECT 127.535 105.945 129.835 106.265 ;
        RECT 150.870 106.385 153.075 106.590 ;
        RECT 127.535 105.425 129.695 105.945 ;
        RECT 150.870 105.930 152.980 106.385 ;
        RECT 8.010 104.590 10.260 104.795 ;
        RECT 19.570 104.740 19.870 105.040 ;
        RECT 21.370 104.740 21.670 105.040 ;
        RECT 21.970 104.740 22.270 105.040 ;
        RECT 22.570 104.740 22.870 105.040 ;
        RECT 23.170 104.740 23.470 105.040 ;
        RECT 24.970 104.740 25.270 105.040 ;
        RECT 8.130 103.905 10.260 104.590 ;
        RECT 21.370 104.140 23.470 104.740 ;
        RECT 31.345 104.590 33.515 105.105 ;
        RECT 31.345 104.265 33.700 104.590 ;
        RECT 8.130 103.690 10.400 103.905 ;
        RECT 21.070 103.840 21.970 104.140 ;
        RECT 22.870 103.840 24.070 104.140 ;
        RECT 8.260 103.010 10.400 103.690 ;
        RECT 20.470 103.540 22.270 103.840 ;
        RECT 22.570 103.540 24.070 103.840 ;
        RECT 31.515 103.760 33.700 104.265 ;
        RECT 20.470 103.240 21.070 103.540 ;
        RECT 21.670 103.240 23.170 103.540 ;
        RECT 23.770 103.240 24.370 103.540 ;
        RECT 31.515 103.425 33.900 103.760 ;
        RECT 8.260 102.795 10.555 103.010 ;
        RECT 20.470 102.940 20.770 103.240 ;
        RECT 8.400 102.120 10.555 102.795 ;
        RECT 20.170 102.640 20.770 102.940 ;
        RECT 20.170 102.340 21.070 102.640 ;
        RECT 21.970 102.340 22.870 103.240 ;
        RECT 24.070 102.940 24.370 103.240 ;
        RECT 24.070 102.640 24.670 102.940 ;
        RECT 23.770 102.340 24.670 102.640 ;
        RECT 31.700 102.930 33.900 103.425 ;
        RECT 31.700 102.590 34.110 102.930 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 127.365 105.105 129.695 105.425 ;
        RECT 139.550 105.485 152.980 105.930 ;
        RECT 139.550 105.480 152.870 105.485 ;
        RECT 127.365 104.590 129.535 105.105 ;
        RECT 127.180 104.265 129.535 104.590 ;
        RECT 135.120 104.700 137.520 105.000 ;
        RECT 135.120 104.400 137.820 104.700 ;
        RECT 127.180 103.760 129.365 104.265 ;
        RECT 134.520 103.800 138.420 104.400 ;
        RECT 139.550 103.930 140.000 105.480 ;
        RECT 150.750 104.795 152.870 105.480 ;
        RECT 150.620 104.590 152.870 104.795 ;
        RECT 150.620 103.905 152.750 104.590 ;
        RECT 126.980 103.425 129.365 103.760 ;
        RECT 126.980 102.930 129.180 103.425 ;
        RECT 8.400 101.905 10.720 102.120 ;
        RECT 8.555 101.235 10.720 101.905 ;
        RECT 8.555 101.010 10.895 101.235 ;
        RECT 20.170 101.140 24.670 102.340 ;
        RECT 31.900 102.105 34.110 102.590 ;
        RECT 31.900 101.760 34.340 102.105 ;
        RECT 32.110 101.285 34.340 101.760 ;
        RECT 8.720 100.350 10.895 101.010 ;
        RECT 8.720 100.120 11.080 100.350 ;
        RECT 8.895 99.465 11.080 100.120 ;
        RECT 18.890 99.550 19.450 100.940 ;
        RECT 20.470 100.540 24.370 101.140 ;
        RECT 32.110 100.930 34.585 101.285 ;
        RECT 21.070 100.240 23.770 100.540 ;
        RECT 21.370 99.940 23.770 100.240 ;
        RECT 32.340 100.470 34.585 100.930 ;
        RECT 32.340 100.105 34.840 100.470 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 126.770 102.590 129.180 102.930 ;
        RECT 134.220 102.600 138.720 103.800 ;
        RECT 150.480 103.690 152.750 103.905 ;
        RECT 150.480 103.010 152.620 103.690 ;
        RECT 126.770 102.105 128.980 102.590 ;
        RECT 126.540 101.760 128.980 102.105 ;
        RECT 134.220 102.300 135.120 102.600 ;
        RECT 134.220 102.000 134.820 102.300 ;
        RECT 126.540 101.285 128.770 101.760 ;
        RECT 134.520 101.700 134.820 102.000 ;
        RECT 136.020 101.700 136.920 102.600 ;
        RECT 137.820 102.300 138.720 102.600 ;
        RECT 138.120 102.000 138.720 102.300 ;
        RECT 150.325 102.795 152.620 103.010 ;
        RECT 150.325 102.120 152.480 102.795 ;
        RECT 138.120 101.700 138.420 102.000 ;
        RECT 134.520 101.400 135.120 101.700 ;
        RECT 135.720 101.400 137.220 101.700 ;
        RECT 137.820 101.400 138.420 101.700 ;
        RECT 126.295 100.930 128.770 101.285 ;
        RECT 134.820 101.100 136.320 101.400 ;
        RECT 136.620 101.100 138.420 101.400 ;
        RECT 150.160 101.905 152.480 102.120 ;
        RECT 150.160 101.235 152.325 101.905 ;
        RECT 126.295 100.470 128.540 100.930 ;
        RECT 134.820 100.800 136.020 101.100 ;
        RECT 136.920 100.800 137.820 101.100 ;
        RECT 149.985 101.010 152.325 101.235 ;
        RECT 32.585 99.660 34.840 100.105 ;
        RECT 8.895 99.235 11.275 99.465 ;
        RECT 9.080 98.585 11.275 99.235 ;
        RECT 18.890 99.120 19.340 99.550 ;
        RECT 32.585 99.285 35.110 99.660 ;
        RECT 32.840 99.120 35.110 99.285 ;
        RECT 18.890 98.855 35.110 99.120 ;
        RECT 18.890 98.670 35.400 98.855 ;
        RECT 9.080 98.350 11.485 98.585 ;
        RECT 32.840 98.470 35.400 98.670 ;
        RECT 9.275 97.705 11.485 98.350 ;
        RECT 33.110 98.050 35.400 98.470 ;
        RECT 9.275 97.580 11.705 97.705 ;
        RECT 33.110 97.660 35.695 98.050 ;
        RECT 9.275 97.465 28.620 97.580 ;
        RECT 9.485 97.130 28.620 97.465 ;
        RECT 9.485 96.830 11.705 97.130 ;
        RECT 9.485 96.585 11.935 96.830 ;
        RECT 9.705 95.960 11.935 96.585 ;
        RECT 23.740 96.350 26.140 96.650 ;
        RECT 23.740 96.050 26.440 96.350 ;
        RECT 9.705 95.705 12.175 95.960 ;
        RECT 9.935 95.090 12.175 95.705 ;
        RECT 23.140 95.450 27.040 96.050 ;
        RECT 28.170 95.580 28.620 97.130 ;
        RECT 33.400 97.255 35.695 97.660 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
        RECT 126.040 100.105 128.540 100.470 ;
        RECT 135.420 100.200 137.520 100.800 ;
        RECT 149.985 100.350 152.160 101.010 ;
        RECT 126.040 99.660 128.295 100.105 ;
        RECT 133.620 99.900 134.520 100.200 ;
        RECT 135.420 99.900 135.720 100.200 ;
        RECT 136.020 99.900 136.320 100.200 ;
        RECT 136.620 99.900 136.920 100.200 ;
        RECT 137.220 99.900 137.520 100.200 ;
        RECT 138.420 99.900 139.320 100.200 ;
        RECT 149.800 100.120 152.160 100.350 ;
        RECT 125.770 99.285 128.295 99.660 ;
        RECT 133.320 99.300 134.820 99.900 ;
        RECT 138.120 99.300 139.620 99.900 ;
        RECT 149.800 99.465 151.985 100.120 ;
        RECT 125.770 98.855 128.040 99.285 ;
        RECT 133.620 99.000 135.420 99.300 ;
        RECT 137.520 99.000 139.320 99.300 ;
        RECT 149.605 99.235 151.985 99.465 ;
        RECT 125.480 98.470 128.040 98.855 ;
        RECT 134.520 98.700 135.720 99.000 ;
        RECT 137.220 98.700 138.420 99.000 ;
        RECT 125.480 98.050 127.770 98.470 ;
        RECT 135.120 98.400 136.320 98.700 ;
        RECT 136.620 98.400 137.820 98.700 ;
        RECT 149.605 98.585 151.800 99.235 ;
        RECT 125.185 97.660 127.770 98.050 ;
        RECT 135.720 97.800 137.220 98.400 ;
        RECT 149.395 98.350 151.800 98.585 ;
        RECT 33.400 96.855 36.010 97.255 ;
        RECT 33.695 96.465 36.010 96.855 ;
        RECT 33.695 96.050 36.340 96.465 ;
        RECT 34.010 95.680 36.340 96.050 ;
        RECT 9.935 94.830 12.430 95.090 ;
        RECT 10.175 94.225 12.430 94.830 ;
        RECT 22.840 94.250 27.340 95.450 ;
        RECT 34.010 95.255 36.680 95.680 ;
        RECT 34.340 94.905 36.680 95.255 ;
        RECT 34.340 94.465 37.035 94.905 ;
        RECT 10.175 93.960 12.690 94.225 ;
        RECT 10.430 93.365 12.690 93.960 ;
        RECT 22.840 93.950 23.740 94.250 ;
        RECT 22.840 93.650 23.440 93.950 ;
        RECT 10.430 93.090 12.965 93.365 ;
        RECT 10.690 92.505 12.965 93.090 ;
        RECT 23.140 93.350 23.440 93.650 ;
        RECT 24.640 93.350 25.540 94.250 ;
        RECT 26.440 93.950 27.340 94.250 ;
        RECT 26.740 93.650 27.340 93.950 ;
        RECT 34.680 94.130 37.035 94.465 ;
        RECT 34.680 93.680 37.400 94.130 ;
        RECT 26.740 93.350 27.040 93.650 ;
        RECT 23.140 93.050 23.740 93.350 ;
        RECT 24.340 93.050 25.840 93.350 ;
        RECT 26.440 93.050 27.040 93.350 ;
        RECT 23.440 92.750 24.940 93.050 ;
        RECT 25.240 92.750 27.040 93.050 ;
        RECT 35.035 93.365 37.400 93.680 ;
        RECT 35.035 92.905 37.785 93.365 ;
        RECT 10.690 92.225 13.250 92.505 ;
        RECT 23.440 92.450 24.640 92.750 ;
        RECT 25.540 92.450 26.440 92.750 ;
        RECT 35.400 92.610 37.785 92.905 ;
        RECT 10.965 91.650 13.250 92.225 ;
        RECT 24.040 91.850 26.140 92.450 ;
        RECT 35.400 92.130 38.180 92.610 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 125.185 97.255 127.480 97.660 ;
        RECT 135.120 97.500 136.320 97.800 ;
        RECT 136.620 97.500 137.820 97.800 ;
        RECT 149.395 97.705 151.605 98.350 ;
        RECT 124.870 96.855 127.480 97.255 ;
        RECT 133.320 97.200 135.720 97.500 ;
        RECT 137.220 97.200 139.320 97.500 ;
        RECT 149.175 97.465 151.605 97.705 ;
        RECT 133.320 96.900 135.120 97.200 ;
        RECT 137.820 96.900 139.620 97.200 ;
        RECT 124.870 96.465 127.185 96.855 ;
        RECT 124.540 96.050 127.185 96.465 ;
        RECT 133.320 96.600 134.520 96.900 ;
        RECT 138.420 96.600 139.620 96.900 ;
        RECT 149.175 96.830 151.395 97.465 ;
        RECT 133.320 96.300 134.220 96.600 ;
        RECT 138.720 96.300 139.620 96.600 ;
        RECT 148.945 96.585 151.395 96.830 ;
        RECT 124.540 95.680 126.870 96.050 ;
        RECT 133.620 96.000 133.920 96.300 ;
        RECT 135.420 96.000 135.720 96.300 ;
        RECT 136.020 96.000 136.320 96.300 ;
        RECT 136.620 96.000 136.920 96.300 ;
        RECT 137.220 96.000 137.520 96.300 ;
        RECT 139.020 96.000 139.320 96.300 ;
        RECT 124.200 95.255 126.870 95.680 ;
        RECT 135.420 95.400 137.520 96.000 ;
        RECT 148.945 95.960 151.175 96.585 ;
        RECT 148.705 95.705 151.175 95.960 ;
        RECT 124.200 94.905 126.540 95.255 ;
        RECT 123.845 94.465 126.540 94.905 ;
        RECT 134.820 95.100 136.020 95.400 ;
        RECT 136.920 95.100 137.820 95.400 ;
        RECT 134.820 94.800 136.320 95.100 ;
        RECT 136.620 94.800 138.420 95.100 ;
        RECT 148.705 95.090 150.945 95.705 ;
        RECT 134.520 94.500 135.120 94.800 ;
        RECT 135.720 94.500 137.220 94.800 ;
        RECT 137.820 94.500 138.420 94.800 ;
        RECT 123.845 94.130 126.200 94.465 ;
        RECT 134.520 94.200 134.820 94.500 ;
        RECT 123.480 93.680 126.200 94.130 ;
        RECT 134.220 93.900 134.820 94.200 ;
        RECT 123.480 93.365 125.845 93.680 ;
        RECT 123.095 92.905 125.845 93.365 ;
        RECT 134.220 93.600 135.120 93.900 ;
        RECT 136.020 93.600 136.920 94.500 ;
        RECT 138.120 94.200 138.420 94.500 ;
        RECT 148.450 94.830 150.945 95.090 ;
        RECT 148.450 94.225 150.705 94.830 ;
        RECT 138.120 93.900 138.720 94.200 ;
        RECT 137.820 93.600 138.720 93.900 ;
        RECT 123.095 92.610 125.480 92.905 ;
        RECT 35.785 91.855 38.180 92.130 ;
        RECT 10.965 91.365 13.545 91.650 ;
        RECT 22.240 91.550 23.140 91.850 ;
        RECT 24.040 91.550 24.340 91.850 ;
        RECT 24.640 91.550 24.940 91.850 ;
        RECT 25.240 91.550 25.540 91.850 ;
        RECT 25.840 91.550 26.140 91.850 ;
        RECT 27.040 91.550 27.940 91.850 ;
        RECT 11.250 90.800 13.545 91.365 ;
        RECT 21.940 90.950 23.440 91.550 ;
        RECT 26.740 90.950 28.240 91.550 ;
        RECT 35.785 91.365 38.585 91.855 ;
        RECT 36.180 91.110 38.585 91.365 ;
        RECT 11.250 90.505 13.855 90.800 ;
        RECT 22.240 90.650 24.040 90.950 ;
        RECT 26.140 90.650 27.940 90.950 ;
        RECT 11.545 89.950 13.855 90.505 ;
        RECT 23.140 90.350 24.340 90.650 ;
        RECT 25.840 90.350 27.040 90.650 ;
        RECT 36.180 90.610 39.005 91.110 ;
        RECT 36.585 90.375 39.005 90.610 ;
        RECT 23.740 90.050 24.940 90.350 ;
        RECT 25.240 90.050 26.440 90.350 ;
        RECT 11.545 89.650 14.170 89.950 ;
        RECT 11.855 89.110 14.170 89.650 ;
        RECT 24.340 89.450 25.840 90.050 ;
        RECT 36.585 89.855 39.440 90.375 ;
        RECT 37.005 89.645 39.440 89.855 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
        RECT 122.700 92.130 125.480 92.610 ;
        RECT 134.220 92.400 138.720 93.600 ;
        RECT 148.190 93.960 150.705 94.225 ;
        RECT 148.190 93.365 150.450 93.960 ;
        RECT 147.915 93.090 150.450 93.365 ;
        RECT 147.915 92.505 150.190 93.090 ;
        RECT 122.700 91.855 125.095 92.130 ;
        RECT 122.295 91.365 125.095 91.855 ;
        RECT 134.520 91.800 138.420 92.400 ;
        RECT 147.630 92.225 150.190 92.505 ;
        RECT 135.120 91.500 137.820 91.800 ;
        RECT 122.295 91.110 124.700 91.365 ;
        RECT 135.120 91.200 137.520 91.500 ;
        RECT 121.875 90.610 124.700 91.110 ;
        RECT 139.440 90.810 140.000 92.200 ;
        RECT 147.630 91.650 149.915 92.225 ;
        RECT 121.875 90.380 124.295 90.610 ;
        RECT 139.550 90.380 140.000 90.810 ;
        RECT 147.335 91.365 149.915 91.650 ;
        RECT 147.335 90.800 149.630 91.365 ;
        RECT 121.875 90.375 140.000 90.380 ;
        RECT 121.440 89.930 140.000 90.375 ;
        RECT 147.025 90.505 149.630 90.800 ;
        RECT 147.025 89.950 149.335 90.505 ;
        RECT 121.440 89.855 124.295 89.930 ;
        RECT 23.740 89.150 24.940 89.450 ;
        RECT 25.240 89.150 26.440 89.450 ;
        RECT 11.855 88.800 14.500 89.110 ;
        RECT 12.170 88.270 14.500 88.800 ;
        RECT 21.940 88.850 24.340 89.150 ;
        RECT 25.840 88.850 27.940 89.150 ;
        RECT 37.005 89.110 39.890 89.645 ;
        RECT 37.440 88.925 39.890 89.110 ;
        RECT 21.940 88.550 23.740 88.850 ;
        RECT 26.440 88.550 28.240 88.850 ;
        RECT 12.170 87.950 14.835 88.270 ;
        RECT 21.940 88.250 23.140 88.550 ;
        RECT 27.040 88.250 28.240 88.550 ;
        RECT 37.440 88.375 40.350 88.925 ;
        RECT 21.940 87.950 22.840 88.250 ;
        RECT 27.340 87.950 28.240 88.250 ;
        RECT 37.890 88.210 40.350 88.375 ;
        RECT 12.500 87.435 14.835 87.950 ;
        RECT 22.240 87.650 22.540 87.950 ;
        RECT 24.040 87.650 24.340 87.950 ;
        RECT 24.640 87.650 24.940 87.950 ;
        RECT 25.240 87.650 25.540 87.950 ;
        RECT 25.840 87.650 26.140 87.950 ;
        RECT 27.640 87.650 27.940 87.950 ;
        RECT 12.500 87.110 15.185 87.435 ;
        RECT 12.835 86.605 15.185 87.110 ;
        RECT 24.040 87.050 26.140 87.650 ;
        RECT 37.890 87.645 40.820 88.210 ;
        RECT 38.350 87.505 40.820 87.645 ;
        RECT 23.440 86.750 24.640 87.050 ;
        RECT 25.540 86.750 26.440 87.050 ;
        RECT 38.350 86.925 41.305 87.505 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 121.440 89.645 123.875 89.855 ;
        RECT 120.990 89.110 123.875 89.645 ;
        RECT 146.710 89.650 149.335 89.950 ;
        RECT 146.710 89.535 149.025 89.650 ;
        RECT 120.990 88.925 123.440 89.110 ;
        RECT 120.530 88.375 123.440 88.925 ;
        RECT 131.790 89.085 149.025 89.535 ;
        RECT 127.360 88.590 129.760 88.890 ;
        RECT 120.530 88.210 122.990 88.375 ;
        RECT 127.360 88.290 130.060 88.590 ;
        RECT 120.060 87.645 122.990 88.210 ;
        RECT 126.760 87.690 130.660 88.290 ;
        RECT 131.790 87.820 132.240 89.085 ;
        RECT 146.380 88.800 149.025 89.085 ;
        RECT 146.380 88.270 148.710 88.800 ;
        RECT 146.045 87.950 148.710 88.270 ;
        RECT 120.060 87.505 122.530 87.645 ;
        RECT 38.820 86.810 41.305 86.925 ;
        RECT 12.835 86.270 15.545 86.605 ;
        RECT 23.440 86.450 24.940 86.750 ;
        RECT 25.240 86.450 27.040 86.750 ;
        RECT 13.185 85.775 15.545 86.270 ;
        RECT 23.140 86.150 23.740 86.450 ;
        RECT 24.340 86.150 25.840 86.450 ;
        RECT 26.440 86.150 27.040 86.450 ;
        RECT 38.820 86.210 41.800 86.810 ;
        RECT 23.140 85.850 23.440 86.150 ;
        RECT 13.185 85.435 15.915 85.775 ;
        RECT 13.545 84.955 15.915 85.435 ;
        RECT 22.840 85.550 23.440 85.850 ;
        RECT 22.840 85.250 23.740 85.550 ;
        RECT 24.640 85.250 25.540 86.150 ;
        RECT 26.740 85.850 27.040 86.150 ;
        RECT 39.305 86.125 41.800 86.210 ;
        RECT 26.740 85.550 27.340 85.850 ;
        RECT 26.440 85.250 27.340 85.550 ;
        RECT 39.305 85.505 42.310 86.125 ;
        RECT 13.545 84.605 16.295 84.955 ;
        RECT 13.915 84.140 16.295 84.605 ;
        RECT 13.915 83.775 16.685 84.140 ;
        RECT 22.840 84.050 27.340 85.250 ;
        RECT 39.800 85.445 42.310 85.505 ;
        RECT 39.800 84.810 42.830 85.445 ;
        RECT 40.310 84.775 42.830 84.810 ;
        RECT 40.310 84.125 43.360 84.775 ;
        RECT 40.830 84.115 43.360 84.125 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 119.575 86.925 122.530 87.505 ;
        RECT 119.575 86.810 122.060 86.925 ;
        RECT 119.080 86.210 122.060 86.810 ;
        RECT 126.460 86.490 130.960 87.690 ;
        RECT 146.045 87.435 148.380 87.950 ;
        RECT 145.695 87.110 148.380 87.435 ;
        RECT 145.695 86.605 148.045 87.110 ;
        RECT 119.080 86.125 121.575 86.210 ;
        RECT 118.570 85.505 121.575 86.125 ;
        RECT 126.460 86.190 127.360 86.490 ;
        RECT 126.460 85.890 127.060 86.190 ;
        RECT 126.760 85.590 127.060 85.890 ;
        RECT 128.260 85.590 129.160 86.490 ;
        RECT 130.060 86.190 130.960 86.490 ;
        RECT 130.360 85.890 130.960 86.190 ;
        RECT 145.335 86.270 148.045 86.605 ;
        RECT 130.360 85.590 130.660 85.890 ;
        RECT 145.335 85.775 147.695 86.270 ;
        RECT 118.570 85.445 121.080 85.505 ;
        RECT 118.050 84.810 121.080 85.445 ;
        RECT 126.760 85.290 127.360 85.590 ;
        RECT 127.960 85.290 129.460 85.590 ;
        RECT 130.060 85.290 130.660 85.590 ;
        RECT 127.060 84.990 128.560 85.290 ;
        RECT 128.860 84.990 130.660 85.290 ;
        RECT 144.965 85.435 147.695 85.775 ;
        RECT 118.050 84.775 120.570 84.810 ;
        RECT 14.295 83.330 16.685 83.775 ;
        RECT 23.140 83.450 27.040 84.050 ;
        RECT 14.295 82.955 17.085 83.330 ;
        RECT 14.685 82.525 17.085 82.955 ;
        RECT 23.740 83.150 26.440 83.450 ;
        RECT 23.740 82.850 26.140 83.150 ;
        RECT 14.685 82.140 17.495 82.525 ;
        RECT 28.060 82.460 28.620 83.850 ;
        RECT 40.830 83.465 43.905 84.115 ;
        RECT 40.830 83.445 44.460 83.465 ;
        RECT 15.085 81.720 17.495 82.140 ;
        RECT 28.170 82.030 28.620 82.460 ;
        RECT 41.235 82.825 44.460 83.445 ;
        RECT 41.235 82.775 45.030 82.825 ;
        RECT 41.235 82.030 41.685 82.775 ;
        RECT 41.905 82.195 45.030 82.775 ;
        RECT 41.905 82.115 45.605 82.195 ;
        RECT 15.085 81.330 17.920 81.720 ;
        RECT 28.170 81.580 41.685 82.030 ;
        RECT 42.460 81.575 45.605 82.115 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
        RECT 117.520 84.125 120.570 84.775 ;
        RECT 127.060 84.690 128.260 84.990 ;
        RECT 129.160 84.690 130.060 84.990 ;
        RECT 144.965 84.955 147.335 85.435 ;
        RECT 117.520 84.115 120.050 84.125 ;
        RECT 116.975 83.465 120.050 84.115 ;
        RECT 127.660 84.090 129.760 84.690 ;
        RECT 144.585 84.605 147.335 84.955 ;
        RECT 144.585 84.140 146.965 84.605 ;
        RECT 125.860 83.790 126.760 84.090 ;
        RECT 127.660 83.790 127.960 84.090 ;
        RECT 128.260 83.790 128.560 84.090 ;
        RECT 128.860 83.790 129.160 84.090 ;
        RECT 129.460 83.790 129.760 84.090 ;
        RECT 130.660 83.790 131.560 84.090 ;
        RECT 116.420 83.445 120.050 83.465 ;
        RECT 116.420 82.825 119.520 83.445 ;
        RECT 125.560 83.190 127.060 83.790 ;
        RECT 130.360 83.190 131.860 83.790 ;
        RECT 144.195 83.775 146.965 84.140 ;
        RECT 144.195 83.330 146.585 83.775 ;
        RECT 125.860 82.890 127.660 83.190 ;
        RECT 129.760 82.890 131.560 83.190 ;
        RECT 143.795 82.955 146.585 83.330 ;
        RECT 115.850 82.775 119.520 82.825 ;
        RECT 115.850 82.195 118.975 82.775 ;
        RECT 126.760 82.590 127.960 82.890 ;
        RECT 129.460 82.590 130.660 82.890 ;
        RECT 127.360 82.290 128.560 82.590 ;
        RECT 128.860 82.290 130.060 82.590 ;
        RECT 143.795 82.525 146.195 82.955 ;
        RECT 42.460 81.465 46.195 81.575 ;
        RECT 15.495 80.925 17.920 81.330 ;
        RECT 43.030 81.245 46.195 81.465 ;
        RECT 38.240 80.965 46.195 81.245 ;
        RECT 15.495 80.525 18.350 80.925 ;
        RECT 15.920 80.135 18.350 80.525 ;
        RECT 38.240 80.795 46.795 80.965 ;
        RECT 15.920 79.720 18.790 80.135 ;
        RECT 38.240 79.920 38.690 80.795 ;
        RECT 43.605 80.365 46.795 80.795 ;
        RECT 43.605 80.195 47.405 80.365 ;
        RECT 16.350 79.350 18.790 79.720 ;
        RECT 16.350 78.925 19.240 79.350 ;
        RECT 33.810 79.230 36.210 79.530 ;
        RECT 33.810 78.930 36.510 79.230 ;
        RECT 16.790 78.575 19.240 78.925 ;
        RECT 16.790 78.135 19.700 78.575 ;
        RECT 33.210 78.330 37.110 78.930 ;
        RECT 38.130 78.530 38.690 79.920 ;
        RECT 44.195 79.775 47.405 80.195 ;
        RECT 44.195 79.575 48.025 79.775 ;
        RECT 44.795 79.200 48.025 79.575 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 115.275 82.115 118.975 82.195 ;
        RECT 115.275 81.575 118.420 82.115 ;
        RECT 127.960 81.690 129.460 82.290 ;
        RECT 143.385 82.140 146.195 82.525 ;
        RECT 143.385 81.720 145.795 82.140 ;
        RECT 114.685 81.465 118.420 81.575 ;
        RECT 114.685 80.965 117.850 81.465 ;
        RECT 127.360 81.390 128.560 81.690 ;
        RECT 128.860 81.390 130.060 81.690 ;
        RECT 114.085 80.825 117.850 80.965 ;
        RECT 125.560 81.090 127.960 81.390 ;
        RECT 129.460 81.090 131.560 81.390 ;
        RECT 142.960 81.330 145.795 81.720 ;
        RECT 114.085 80.365 117.275 80.825 ;
        RECT 113.475 80.195 117.275 80.365 ;
        RECT 125.560 80.790 127.360 81.090 ;
        RECT 130.060 80.790 131.860 81.090 ;
        RECT 142.960 80.925 145.385 81.330 ;
        RECT 125.560 80.490 126.760 80.790 ;
        RECT 130.660 80.490 131.860 80.790 ;
        RECT 113.475 79.775 116.685 80.195 ;
        RECT 125.560 80.190 126.460 80.490 ;
        RECT 130.960 80.190 131.860 80.490 ;
        RECT 142.530 80.525 145.385 80.925 ;
        RECT 125.860 79.890 126.160 80.190 ;
        RECT 127.660 79.890 127.960 80.190 ;
        RECT 128.260 79.890 128.560 80.190 ;
        RECT 128.860 79.890 129.160 80.190 ;
        RECT 129.460 79.890 129.760 80.190 ;
        RECT 131.260 79.890 131.560 80.190 ;
        RECT 142.530 80.135 144.960 80.525 ;
        RECT 112.855 79.575 116.685 79.775 ;
        RECT 44.795 78.965 48.655 79.200 ;
        RECT 45.405 78.630 48.655 78.965 ;
        RECT 45.405 78.365 49.295 78.630 ;
        RECT 17.240 77.800 19.700 78.135 ;
        RECT 17.240 77.350 20.170 77.800 ;
        RECT 17.700 77.035 20.170 77.350 ;
        RECT 32.910 77.130 37.410 78.330 ;
        RECT 46.025 78.075 49.295 78.365 ;
        RECT 46.025 77.775 49.945 78.075 ;
        RECT 46.655 77.530 49.945 77.775 ;
        RECT 46.655 77.200 50.605 77.530 ;
        RECT 17.700 76.575 20.650 77.035 ;
        RECT 18.170 76.270 20.650 76.575 ;
        RECT 32.910 76.830 33.810 77.130 ;
        RECT 32.910 76.530 33.510 76.830 ;
        RECT 18.170 75.800 21.140 76.270 ;
        RECT 33.210 76.230 33.510 76.530 ;
        RECT 34.710 76.230 35.610 77.130 ;
        RECT 36.510 76.830 37.410 77.130 ;
        RECT 36.810 76.530 37.410 76.830 ;
        RECT 47.295 77.000 50.605 77.200 ;
        RECT 47.295 76.630 51.275 77.000 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
        RECT 112.855 79.200 116.085 79.575 ;
        RECT 127.660 79.290 129.760 79.890 ;
        RECT 142.090 79.720 144.960 80.135 ;
        RECT 142.090 79.350 144.530 79.720 ;
        RECT 112.225 78.965 116.085 79.200 ;
        RECT 127.060 78.990 128.260 79.290 ;
        RECT 129.160 78.990 130.060 79.290 ;
        RECT 112.225 78.630 115.475 78.965 ;
        RECT 127.060 78.690 128.560 78.990 ;
        RECT 128.860 78.690 130.660 78.990 ;
        RECT 111.585 78.365 115.475 78.630 ;
        RECT 126.760 78.390 127.360 78.690 ;
        RECT 127.960 78.390 129.460 78.690 ;
        RECT 130.060 78.390 130.660 78.690 ;
        RECT 141.640 78.925 144.530 79.350 ;
        RECT 141.640 78.575 144.090 78.925 ;
        RECT 111.585 78.075 114.855 78.365 ;
        RECT 126.760 78.090 127.060 78.390 ;
        RECT 110.935 77.775 114.855 78.075 ;
        RECT 126.460 77.790 127.060 78.090 ;
        RECT 110.935 77.530 114.225 77.775 ;
        RECT 110.275 77.200 114.225 77.530 ;
        RECT 126.460 77.490 127.360 77.790 ;
        RECT 128.260 77.490 129.160 78.390 ;
        RECT 130.360 78.090 130.660 78.390 ;
        RECT 141.180 78.135 144.090 78.575 ;
        RECT 130.360 77.790 130.960 78.090 ;
        RECT 141.180 77.800 143.640 78.135 ;
        RECT 130.060 77.490 130.960 77.790 ;
        RECT 110.275 77.000 113.585 77.200 ;
        RECT 36.810 76.230 37.110 76.530 ;
        RECT 33.210 75.930 33.810 76.230 ;
        RECT 34.410 75.930 35.910 76.230 ;
        RECT 36.510 75.930 37.110 76.230 ;
        RECT 47.945 76.480 51.275 76.630 ;
        RECT 109.605 76.630 113.585 77.000 ;
        RECT 109.605 76.480 112.935 76.630 ;
        RECT 47.945 76.075 51.955 76.480 ;
        RECT 18.650 75.515 21.140 75.800 ;
        RECT 33.510 75.630 35.010 75.930 ;
        RECT 35.310 75.630 37.110 75.930 ;
        RECT 48.605 75.970 51.955 76.075 ;
        RECT 108.925 76.075 112.935 76.480 ;
        RECT 126.460 76.290 130.960 77.490 ;
        RECT 140.710 77.350 143.640 77.800 ;
        RECT 140.710 77.035 143.180 77.350 ;
        RECT 140.230 76.575 143.180 77.035 ;
        RECT 108.925 75.970 112.275 76.075 ;
        RECT 18.650 75.035 21.640 75.515 ;
        RECT 33.510 75.330 34.710 75.630 ;
        RECT 35.610 75.330 36.510 75.630 ;
        RECT 48.605 75.530 52.640 75.970 ;
        RECT 49.275 75.475 52.640 75.530 ;
        RECT 108.240 75.530 112.275 75.970 ;
        RECT 126.760 75.690 130.660 76.290 ;
        RECT 140.230 76.270 142.710 76.575 ;
        RECT 108.240 75.475 111.605 75.530 ;
        RECT 19.140 74.770 21.640 75.035 ;
        RECT 19.140 74.270 22.150 74.770 ;
        RECT 34.110 74.730 36.210 75.330 ;
        RECT 49.275 75.000 53.335 75.475 ;
        RECT 49.955 74.990 53.335 75.000 ;
        RECT 107.545 75.000 111.605 75.475 ;
        RECT 127.360 75.390 130.060 75.690 ;
        RECT 127.360 75.090 129.760 75.390 ;
        RECT 107.545 74.990 110.925 75.000 ;
        RECT 32.310 74.430 32.610 74.730 ;
        RECT 34.110 74.430 34.410 74.730 ;
        RECT 34.710 74.430 35.010 74.730 ;
        RECT 35.310 74.430 35.610 74.730 ;
        RECT 35.910 74.430 36.210 74.730 ;
        RECT 37.710 74.430 38.010 74.730 ;
        RECT 49.955 74.520 54.040 74.990 ;
        RECT 106.840 74.520 110.925 74.990 ;
        RECT 131.680 74.700 132.240 76.090 ;
        RECT 139.740 75.800 142.710 76.270 ;
        RECT 139.740 75.515 142.230 75.800 ;
        RECT 139.240 75.035 142.230 75.515 ;
        RECT 139.240 74.770 141.740 75.035 ;
        RECT 49.955 74.480 54.755 74.520 ;
        RECT 19.640 74.025 22.150 74.270 ;
        RECT 32.010 74.130 32.910 74.430 ;
        RECT 37.410 74.130 38.310 74.430 ;
        RECT 19.640 73.515 22.665 74.025 ;
        RECT 20.150 73.290 22.665 73.515 ;
        RECT 32.010 73.830 33.210 74.130 ;
        RECT 37.110 73.830 38.310 74.130 ;
        RECT 50.640 74.060 54.755 74.480 ;
        RECT 106.125 74.480 110.925 74.520 ;
        RECT 106.125 74.270 110.240 74.480 ;
        RECT 131.790 74.270 132.240 74.700 ;
        RECT 106.125 74.060 132.240 74.270 ;
        RECT 50.640 73.970 55.475 74.060 ;
        RECT 32.010 73.530 33.810 73.830 ;
        RECT 36.510 73.530 38.310 73.830 ;
        RECT 51.335 73.610 55.475 73.970 ;
        RECT 105.405 73.820 132.240 74.060 ;
        RECT 138.730 74.270 141.740 74.770 ;
        RECT 138.730 74.025 141.240 74.270 ;
        RECT 105.405 73.610 109.545 73.820 ;
        RECT 20.150 72.770 23.195 73.290 ;
        RECT 32.010 73.230 34.410 73.530 ;
        RECT 35.910 73.230 38.010 73.530 ;
        RECT 51.335 73.475 56.205 73.610 ;
        RECT 33.810 72.930 35.010 73.230 ;
        RECT 35.310 72.930 36.510 73.230 ;
        RECT 52.040 73.175 56.205 73.475 ;
        RECT 104.675 73.475 109.545 73.610 ;
        RECT 104.675 73.175 108.840 73.475 ;
        RECT 52.040 72.990 56.940 73.175 ;
        RECT 20.665 72.565 23.195 72.770 ;
        RECT 20.665 72.025 23.730 72.565 ;
        RECT 34.410 72.330 35.910 72.930 ;
        RECT 52.220 72.755 56.940 72.990 ;
        RECT 103.940 72.990 108.840 73.175 ;
        RECT 115.190 73.140 117.590 73.440 ;
        RECT 103.940 72.755 108.125 72.990 ;
        RECT 115.190 72.840 117.890 73.140 ;
        RECT 52.220 72.520 57.685 72.755 ;
        RECT 33.810 72.030 35.010 72.330 ;
        RECT 35.310 72.030 36.510 72.330 ;
        RECT 21.195 71.840 23.730 72.025 ;
        RECT 21.195 71.290 24.275 71.840 ;
        RECT 33.210 71.730 34.410 72.030 ;
        RECT 35.910 71.730 37.110 72.030 ;
        RECT 32.310 71.430 34.110 71.730 ;
        RECT 36.210 71.430 38.010 71.730 ;
        RECT 21.730 71.125 24.275 71.290 ;
        RECT 21.730 70.565 24.830 71.125 ;
        RECT 32.010 70.830 33.510 71.430 ;
        RECT 36.810 70.830 38.310 71.430 ;
        RECT 22.275 70.420 24.830 70.565 ;
        RECT 32.310 70.530 33.210 70.830 ;
        RECT 34.110 70.530 34.410 70.830 ;
        RECT 34.710 70.530 35.010 70.830 ;
        RECT 35.310 70.530 35.610 70.830 ;
        RECT 35.910 70.530 36.210 70.830 ;
        RECT 37.110 70.530 38.010 70.830 ;
        RECT 22.275 69.840 25.395 70.420 ;
        RECT 34.110 69.930 36.210 70.530 ;
        RECT 22.830 69.720 25.395 69.840 ;
        RECT 22.830 69.125 25.965 69.720 ;
        RECT 33.510 69.630 34.710 69.930 ;
        RECT 35.610 69.630 36.510 69.930 ;
        RECT 33.510 69.330 35.010 69.630 ;
        RECT 35.310 69.330 37.110 69.630 ;
        RECT 23.395 69.025 25.965 69.125 ;
        RECT 33.210 69.030 33.810 69.330 ;
        RECT 34.410 69.030 35.910 69.330 ;
        RECT 36.510 69.030 37.110 69.330 ;
        RECT 23.395 68.420 26.545 69.025 ;
        RECT 33.210 68.730 33.510 69.030 ;
        RECT 23.965 68.340 26.545 68.420 ;
        RECT 32.910 68.430 33.510 68.730 ;
        RECT 23.965 67.720 27.135 68.340 ;
        RECT 24.545 67.660 27.135 67.720 ;
        RECT 32.910 68.130 33.810 68.430 ;
        RECT 34.710 68.130 35.610 69.030 ;
        RECT 36.810 68.730 37.110 69.030 ;
        RECT 52.220 68.770 52.670 72.520 ;
        RECT 53.475 72.350 57.685 72.520 ;
        RECT 103.195 72.520 108.125 72.755 ;
        RECT 103.195 72.350 107.405 72.520 ;
        RECT 53.475 72.060 58.440 72.350 ;
        RECT 54.205 71.955 58.440 72.060 ;
        RECT 102.440 72.060 107.405 72.350 ;
        RECT 114.590 72.240 118.490 72.840 ;
        RECT 119.510 72.440 120.070 73.820 ;
        RECT 138.215 73.515 141.240 74.025 ;
        RECT 138.215 73.290 140.730 73.515 ;
        RECT 137.685 72.770 140.730 73.290 ;
        RECT 137.685 72.565 140.215 72.770 ;
        RECT 102.440 71.955 106.675 72.060 ;
        RECT 54.205 71.610 59.195 71.955 ;
        RECT 54.940 71.570 59.195 71.610 ;
        RECT 101.685 71.610 106.675 71.955 ;
        RECT 101.685 71.570 105.940 71.610 ;
        RECT 54.940 71.205 59.960 71.570 ;
        RECT 100.920 71.205 105.940 71.570 ;
        RECT 54.940 71.175 60.735 71.205 ;
        RECT 55.685 70.850 60.735 71.175 ;
        RECT 100.145 71.175 105.940 71.205 ;
        RECT 100.145 70.850 105.195 71.175 ;
        RECT 55.685 70.755 61.510 70.850 ;
        RECT 56.440 70.510 61.510 70.755 ;
        RECT 99.370 70.755 105.195 70.850 ;
        RECT 114.290 71.040 118.790 72.240 ;
        RECT 137.150 72.025 140.215 72.565 ;
        RECT 137.150 71.840 139.685 72.025 ;
        RECT 136.605 71.290 139.685 71.840 ;
        RECT 136.605 71.125 139.150 71.290 ;
        RECT 99.370 70.510 104.590 70.755 ;
        RECT 56.440 70.350 62.295 70.510 ;
        RECT 57.195 70.180 62.295 70.350 ;
        RECT 98.585 70.350 104.590 70.510 ;
        RECT 114.290 70.740 115.190 71.040 ;
        RECT 114.290 70.440 114.890 70.740 ;
        RECT 98.585 70.180 103.685 70.350 ;
        RECT 57.195 69.955 63.085 70.180 ;
        RECT 57.960 69.865 63.085 69.955 ;
        RECT 97.795 69.955 103.685 70.180 ;
        RECT 97.795 69.865 102.920 69.955 ;
        RECT 57.960 69.570 63.880 69.865 ;
        RECT 97.000 69.570 102.920 69.865 ;
        RECT 58.735 69.280 64.685 69.570 ;
        RECT 96.195 69.280 102.145 69.570 ;
        RECT 58.735 69.205 65.490 69.280 ;
        RECT 59.510 69.010 65.490 69.205 ;
        RECT 95.390 69.205 102.145 69.280 ;
        RECT 95.390 69.010 101.370 69.205 ;
        RECT 59.510 68.850 66.300 69.010 ;
        RECT 36.810 68.430 37.410 68.730 ;
        RECT 36.510 68.130 37.410 68.430 ;
        RECT 24.545 67.025 27.735 67.660 ;
        RECT 25.135 66.990 27.735 67.025 ;
        RECT 25.135 66.340 28.340 66.990 ;
        RECT 32.910 66.930 37.410 68.130 ;
        RECT 47.790 68.080 50.190 68.380 ;
        RECT 47.790 67.780 50.490 68.080 ;
        RECT 47.190 67.180 51.090 67.780 ;
        RECT 52.110 67.380 52.670 68.770 ;
        RECT 60.295 68.755 66.300 68.850 ;
        RECT 94.580 68.850 101.370 69.010 ;
        RECT 94.580 68.755 100.585 68.850 ;
        RECT 60.295 68.510 67.115 68.755 ;
        RECT 93.765 68.510 100.585 68.755 ;
        RECT 61.085 68.280 67.935 68.510 ;
        RECT 92.945 68.280 99.795 68.510 ;
        RECT 61.085 68.180 68.760 68.280 ;
        RECT 61.880 68.070 68.760 68.180 ;
        RECT 92.120 68.180 99.795 68.280 ;
        RECT 92.120 68.070 99.000 68.180 ;
        RECT 61.880 67.870 69.590 68.070 ;
        RECT 91.290 67.870 99.000 68.070 ;
        RECT 61.880 67.865 70.420 67.870 ;
        RECT 62.685 67.685 70.420 67.865 ;
        RECT 90.460 67.865 99.000 67.870 ;
        RECT 90.460 67.685 98.195 67.865 ;
        RECT 62.685 67.570 71.255 67.685 ;
        RECT 63.490 67.515 71.255 67.570 ;
        RECT 89.625 67.570 98.195 67.685 ;
        RECT 89.625 67.515 97.390 67.570 ;
        RECT 63.490 67.355 72.095 67.515 ;
        RECT 88.785 67.355 97.390 67.515 ;
        RECT 63.490 67.280 72.935 67.355 ;
        RECT 64.300 67.215 72.935 67.280 ;
        RECT 87.945 67.280 97.390 67.355 ;
        RECT 87.945 67.215 96.580 67.280 ;
        RECT 25.735 66.325 28.340 66.340 ;
        RECT 33.210 66.330 37.110 66.930 ;
        RECT 25.735 65.670 28.955 66.325 ;
        RECT 33.810 66.030 36.510 66.330 ;
        RECT 33.810 65.730 36.210 66.030 ;
        RECT 25.735 65.660 29.580 65.670 ;
        RECT 26.340 65.020 29.580 65.660 ;
        RECT 26.340 64.990 30.210 65.020 ;
        RECT 26.955 64.380 30.210 64.990 ;
        RECT 26.955 64.325 30.850 64.380 ;
        RECT 27.580 63.750 30.850 64.325 ;
        RECT 27.580 63.670 31.500 63.750 ;
        RECT 28.210 63.125 31.500 63.670 ;
        RECT 28.210 63.020 32.155 63.125 ;
        RECT 28.850 62.510 32.155 63.020 ;
        RECT 28.850 62.380 32.820 62.510 ;
        RECT 29.500 61.905 32.820 62.380 ;
        RECT 29.500 61.750 33.490 61.905 ;
        RECT 30.155 61.305 33.490 61.750 ;
        RECT 30.155 61.125 34.170 61.305 ;
        RECT 30.820 60.715 34.170 61.125 ;
        RECT 30.820 60.510 34.855 60.715 ;
        RECT 31.490 60.135 34.855 60.510 ;
        RECT 31.490 59.905 35.550 60.135 ;
        RECT 32.170 59.565 35.550 59.905 ;
        RECT 32.170 59.305 36.250 59.565 ;
        RECT 32.855 59.000 36.250 59.305 ;
        RECT 32.855 58.715 36.955 59.000 ;
        RECT 33.550 58.445 36.955 58.715 ;
        RECT 33.550 58.135 37.670 58.445 ;
        RECT 34.250 57.900 37.670 58.135 ;
        RECT 38.240 57.900 38.690 66.800 ;
        RECT 46.890 65.980 51.390 67.180 ;
        RECT 64.300 67.090 73.775 67.215 ;
        RECT 87.105 67.090 96.580 67.215 ;
        RECT 64.300 67.010 74.625 67.090 ;
        RECT 65.115 66.980 74.625 67.010 ;
        RECT 86.255 67.010 96.580 67.090 ;
        RECT 86.255 66.980 95.765 67.010 ;
        RECT 65.115 66.880 75.470 66.980 ;
        RECT 85.410 66.880 95.765 66.980 ;
        RECT 65.115 66.800 76.320 66.880 ;
        RECT 84.560 66.800 95.765 66.880 ;
        RECT 65.115 66.755 77.170 66.800 ;
        RECT 65.935 66.730 77.170 66.755 ;
        RECT 83.710 66.755 95.765 66.800 ;
        RECT 83.710 66.730 94.945 66.755 ;
        RECT 65.935 66.680 78.025 66.730 ;
        RECT 82.855 66.680 94.945 66.730 ;
        RECT 65.935 66.640 78.880 66.680 ;
        RECT 82.000 66.640 94.945 66.680 ;
        RECT 65.935 66.620 79.730 66.640 ;
        RECT 81.150 66.620 94.945 66.640 ;
        RECT 65.935 66.510 94.945 66.620 ;
        RECT 66.760 66.280 94.120 66.510 ;
        RECT 67.590 66.070 93.290 66.280 ;
        RECT 46.890 65.680 47.790 65.980 ;
        RECT 46.890 65.380 47.490 65.680 ;
        RECT 47.190 65.080 47.490 65.380 ;
        RECT 48.690 65.080 49.590 65.980 ;
        RECT 50.490 65.680 51.390 65.980 ;
        RECT 68.420 65.870 92.460 66.070 ;
        RECT 50.790 65.380 51.390 65.680 ;
        RECT 68.870 65.685 91.625 65.870 ;
        RECT 50.790 65.080 51.090 65.380 ;
        RECT 47.190 64.780 47.790 65.080 ;
        RECT 48.390 64.780 49.890 65.080 ;
        RECT 50.490 64.780 51.090 65.080 ;
        RECT 47.490 64.480 48.990 64.780 ;
        RECT 49.290 64.480 51.090 64.780 ;
        RECT 47.490 64.180 48.690 64.480 ;
        RECT 49.590 64.180 50.490 64.480 ;
        RECT 48.090 63.580 50.190 64.180 ;
        RECT 46.290 63.280 46.590 63.580 ;
        RECT 48.090 63.280 48.390 63.580 ;
        RECT 48.690 63.280 48.990 63.580 ;
        RECT 49.290 63.280 49.590 63.580 ;
        RECT 49.890 63.280 50.190 63.580 ;
        RECT 51.690 63.280 51.990 63.580 ;
        RECT 45.990 62.980 46.890 63.280 ;
        RECT 51.390 62.980 52.290 63.280 ;
        RECT 45.990 62.680 47.190 62.980 ;
        RECT 51.090 62.680 52.290 62.980 ;
        RECT 45.990 62.380 47.790 62.680 ;
        RECT 50.490 62.380 52.290 62.680 ;
        RECT 45.990 62.080 48.390 62.380 ;
        RECT 49.890 62.080 51.990 62.380 ;
        RECT 68.870 62.240 69.320 65.685 ;
        RECT 70.095 65.515 90.785 65.685 ;
        RECT 70.935 65.355 89.945 65.515 ;
        RECT 71.775 65.215 89.105 65.355 ;
        RECT 72.625 65.090 88.255 65.215 ;
        RECT 73.470 64.980 87.410 65.090 ;
        RECT 74.320 64.880 86.560 64.980 ;
        RECT 75.170 64.800 85.710 64.880 ;
        RECT 76.025 64.730 84.855 64.800 ;
        RECT 76.880 64.680 84.000 64.730 ;
        RECT 77.730 64.640 83.150 64.680 ;
        RECT 78.585 64.620 82.295 64.640 ;
        RECT 79.440 64.610 81.435 64.620 ;
        RECT 47.790 61.780 48.990 62.080 ;
        RECT 49.290 61.780 50.490 62.080 ;
        RECT 48.390 61.180 49.890 61.780 ;
        RECT 64.440 61.550 66.840 61.850 ;
        RECT 64.440 61.250 67.140 61.550 ;
        RECT 47.790 60.880 48.990 61.180 ;
        RECT 49.290 60.880 50.490 61.180 ;
        RECT 47.190 60.580 48.390 60.880 ;
        RECT 49.890 60.580 51.090 60.880 ;
        RECT 63.840 60.650 67.740 61.250 ;
        RECT 68.760 60.850 69.320 62.240 ;
        RECT 86.700 60.900 87.150 64.980 ;
        RECT 104.140 64.880 104.590 70.350 ;
        RECT 114.590 70.140 114.890 70.440 ;
        RECT 116.090 70.140 116.990 71.040 ;
        RECT 117.890 70.740 118.790 71.040 ;
        RECT 118.190 70.440 118.790 70.740 ;
        RECT 136.050 70.565 139.150 71.125 ;
        RECT 118.190 70.140 118.490 70.440 ;
        RECT 136.050 70.420 138.605 70.565 ;
        RECT 114.590 69.840 115.190 70.140 ;
        RECT 115.790 69.840 117.290 70.140 ;
        RECT 117.890 69.840 118.490 70.140 ;
        RECT 114.890 69.540 116.390 69.840 ;
        RECT 116.690 69.540 118.490 69.840 ;
        RECT 135.485 69.840 138.605 70.420 ;
        RECT 135.485 69.720 138.050 69.840 ;
        RECT 114.890 69.240 116.090 69.540 ;
        RECT 116.990 69.240 117.890 69.540 ;
        RECT 115.490 68.640 117.590 69.240 ;
        RECT 134.915 69.125 138.050 69.720 ;
        RECT 134.915 69.025 137.485 69.125 ;
        RECT 113.690 68.340 113.990 68.640 ;
        RECT 115.490 68.340 115.790 68.640 ;
        RECT 116.090 68.340 116.390 68.640 ;
        RECT 116.690 68.340 116.990 68.640 ;
        RECT 117.290 68.340 117.590 68.640 ;
        RECT 119.090 68.340 119.390 68.640 ;
        RECT 134.335 68.420 137.485 69.025 ;
        RECT 134.335 68.340 136.915 68.420 ;
        RECT 113.390 68.040 114.290 68.340 ;
        RECT 118.790 68.040 119.690 68.340 ;
        RECT 113.390 67.740 114.590 68.040 ;
        RECT 118.490 67.740 119.690 68.040 ;
        RECT 113.390 67.440 115.190 67.740 ;
        RECT 117.890 67.440 119.690 67.740 ;
        RECT 133.745 67.720 136.915 68.340 ;
        RECT 133.745 67.660 136.335 67.720 ;
        RECT 113.390 67.140 115.790 67.440 ;
        RECT 117.290 67.140 119.390 67.440 ;
        RECT 115.190 66.840 116.390 67.140 ;
        RECT 116.690 66.840 117.890 67.140 ;
        RECT 133.145 67.025 136.335 67.660 ;
        RECT 133.145 66.990 135.745 67.025 ;
        RECT 115.790 66.240 117.290 66.840 ;
        RECT 132.540 66.340 135.745 66.990 ;
        RECT 132.540 66.325 135.145 66.340 ;
        RECT 115.190 65.940 116.390 66.240 ;
        RECT 116.690 65.940 117.890 66.240 ;
        RECT 114.590 65.640 115.790 65.940 ;
        RECT 117.290 65.640 118.490 65.940 ;
        RECT 131.925 65.670 135.145 66.325 ;
        RECT 131.300 65.660 135.145 65.670 ;
        RECT 113.690 65.340 115.490 65.640 ;
        RECT 117.590 65.340 119.390 65.640 ;
        RECT 99.710 64.190 102.110 64.490 ;
        RECT 99.710 63.890 102.410 64.190 ;
        RECT 99.110 63.290 103.010 63.890 ;
        RECT 104.030 63.490 104.590 64.880 ;
        RECT 113.390 64.740 114.890 65.340 ;
        RECT 118.190 64.740 119.690 65.340 ;
        RECT 131.300 65.020 134.540 65.660 ;
        RECT 130.670 64.990 134.540 65.020 ;
        RECT 113.690 64.440 114.590 64.740 ;
        RECT 115.490 64.440 115.790 64.740 ;
        RECT 116.090 64.440 116.390 64.740 ;
        RECT 116.690 64.440 116.990 64.740 ;
        RECT 117.290 64.440 117.590 64.740 ;
        RECT 118.490 64.440 119.390 64.740 ;
        RECT 115.490 63.840 117.590 64.440 ;
        RECT 130.670 64.380 133.925 64.990 ;
        RECT 130.030 64.325 133.925 64.380 ;
        RECT 114.890 63.540 116.090 63.840 ;
        RECT 116.990 63.540 117.890 63.840 ;
        RECT 130.030 63.750 133.300 64.325 ;
        RECT 129.380 63.670 133.300 63.750 ;
        RECT 98.810 62.090 103.310 63.290 ;
        RECT 114.890 63.240 116.390 63.540 ;
        RECT 116.690 63.240 118.490 63.540 ;
        RECT 114.590 62.940 115.190 63.240 ;
        RECT 115.790 62.940 117.290 63.240 ;
        RECT 117.890 62.940 118.490 63.240 ;
        RECT 129.380 63.125 132.670 63.670 ;
        RECT 114.590 62.640 114.890 62.940 ;
        RECT 98.810 61.790 99.710 62.090 ;
        RECT 98.810 61.490 99.410 61.790 ;
        RECT 46.290 60.280 48.090 60.580 ;
        RECT 50.190 60.280 51.990 60.580 ;
        RECT 45.990 59.680 47.490 60.280 ;
        RECT 50.790 59.680 52.290 60.280 ;
        RECT 46.290 59.380 47.190 59.680 ;
        RECT 48.090 59.380 48.390 59.680 ;
        RECT 48.690 59.380 48.990 59.680 ;
        RECT 49.290 59.380 49.590 59.680 ;
        RECT 49.890 59.380 50.190 59.680 ;
        RECT 51.090 59.380 51.990 59.680 ;
        RECT 63.540 59.450 68.040 60.650 ;
        RECT 82.270 60.210 84.670 60.510 ;
        RECT 82.270 59.910 84.970 60.210 ;
        RECT 48.090 58.780 50.190 59.380 ;
        RECT 63.540 59.150 64.440 59.450 ;
        RECT 63.540 58.850 64.140 59.150 ;
        RECT 47.490 58.480 48.690 58.780 ;
        RECT 49.590 58.480 50.490 58.780 ;
        RECT 63.840 58.550 64.140 58.850 ;
        RECT 65.340 58.550 66.240 59.450 ;
        RECT 67.140 59.150 68.040 59.450 ;
        RECT 81.670 59.310 85.570 59.910 ;
        RECT 86.590 59.510 87.150 60.900 ;
        RECT 99.110 61.190 99.410 61.490 ;
        RECT 100.610 61.190 101.510 62.090 ;
        RECT 102.410 61.790 103.310 62.090 ;
        RECT 102.710 61.490 103.310 61.790 ;
        RECT 114.290 62.340 114.890 62.640 ;
        RECT 114.290 62.040 115.190 62.340 ;
        RECT 116.090 62.040 116.990 62.940 ;
        RECT 118.190 62.640 118.490 62.940 ;
        RECT 128.725 63.020 132.670 63.125 ;
        RECT 118.190 62.340 118.790 62.640 ;
        RECT 128.725 62.510 132.030 63.020 ;
        RECT 117.890 62.040 118.790 62.340 ;
        RECT 102.710 61.190 103.010 61.490 ;
        RECT 99.110 60.890 99.710 61.190 ;
        RECT 100.310 60.890 101.810 61.190 ;
        RECT 102.410 60.890 103.010 61.190 ;
        RECT 99.410 60.590 100.910 60.890 ;
        RECT 101.210 60.590 103.010 60.890 ;
        RECT 114.290 60.840 118.790 62.040 ;
        RECT 128.060 62.380 132.030 62.510 ;
        RECT 128.060 61.905 131.380 62.380 ;
        RECT 127.390 61.750 131.380 61.905 ;
        RECT 127.390 61.305 130.725 61.750 ;
        RECT 126.710 61.125 130.725 61.305 ;
        RECT 99.410 60.290 100.610 60.590 ;
        RECT 101.510 60.290 102.410 60.590 ;
        RECT 100.010 59.690 102.110 60.290 ;
        RECT 114.590 60.240 118.490 60.840 ;
        RECT 126.710 60.715 130.060 61.125 ;
        RECT 115.190 59.940 117.890 60.240 ;
        RECT 98.210 59.390 98.510 59.690 ;
        RECT 100.010 59.390 100.310 59.690 ;
        RECT 100.610 59.390 100.910 59.690 ;
        RECT 101.210 59.390 101.510 59.690 ;
        RECT 101.810 59.390 102.110 59.690 ;
        RECT 103.610 59.390 103.910 59.690 ;
        RECT 115.190 59.640 117.590 59.940 ;
        RECT 67.440 58.850 68.040 59.150 ;
        RECT 67.440 58.550 67.740 58.850 ;
        RECT 47.490 58.180 48.990 58.480 ;
        RECT 49.290 58.180 51.090 58.480 ;
        RECT 63.840 58.250 64.440 58.550 ;
        RECT 65.040 58.250 66.540 58.550 ;
        RECT 67.140 58.250 67.740 58.550 ;
        RECT 34.250 57.565 38.690 57.900 ;
        RECT 47.190 57.880 47.790 58.180 ;
        RECT 48.390 57.880 49.890 58.180 ;
        RECT 50.490 57.880 51.090 58.180 ;
        RECT 47.190 57.580 47.490 57.880 ;
        RECT 34.955 57.365 38.690 57.565 ;
        RECT 34.955 57.000 39.120 57.365 ;
        RECT 35.670 56.835 39.120 57.000 ;
        RECT 46.890 57.280 47.490 57.580 ;
        RECT 46.890 56.980 47.790 57.280 ;
        RECT 48.690 56.980 49.590 57.880 ;
        RECT 50.790 57.580 51.090 57.880 ;
        RECT 64.140 57.950 65.640 58.250 ;
        RECT 65.940 57.950 67.740 58.250 ;
        RECT 81.370 58.110 85.870 59.310 ;
        RECT 97.910 59.090 98.810 59.390 ;
        RECT 103.310 59.090 104.210 59.390 ;
        RECT 97.910 58.790 99.110 59.090 ;
        RECT 103.010 58.790 104.210 59.090 ;
        RECT 97.910 58.490 99.710 58.790 ;
        RECT 102.410 58.490 104.210 58.790 ;
        RECT 119.620 59.160 120.070 60.710 ;
        RECT 126.025 60.510 130.060 60.715 ;
        RECT 126.025 60.135 129.390 60.510 ;
        RECT 125.330 59.905 129.390 60.135 ;
        RECT 125.330 59.565 128.710 59.905 ;
        RECT 124.630 59.305 128.710 59.565 ;
        RECT 124.630 59.160 128.025 59.305 ;
        RECT 119.620 58.715 128.025 59.160 ;
        RECT 119.620 58.710 127.330 58.715 ;
        RECT 97.910 58.190 100.310 58.490 ;
        RECT 101.810 58.190 103.910 58.490 ;
        RECT 123.925 58.445 127.330 58.710 ;
        RECT 64.140 57.650 65.340 57.950 ;
        RECT 66.240 57.650 67.140 57.950 ;
        RECT 81.370 57.810 82.270 58.110 ;
        RECT 50.790 57.280 51.390 57.580 ;
        RECT 50.490 56.980 51.390 57.280 ;
        RECT 64.740 57.050 66.840 57.650 ;
        RECT 81.370 57.510 81.970 57.810 ;
        RECT 81.670 57.210 81.970 57.510 ;
        RECT 83.170 57.210 84.070 58.110 ;
        RECT 84.970 57.810 85.870 58.110 ;
        RECT 99.710 57.890 100.910 58.190 ;
        RECT 101.210 57.890 102.410 58.190 ;
        RECT 123.210 58.135 127.330 58.445 ;
        RECT 123.210 57.900 126.630 58.135 ;
        RECT 85.270 57.510 85.870 57.810 ;
        RECT 85.270 57.210 85.570 57.510 ;
        RECT 100.310 57.290 101.810 57.890 ;
        RECT 122.485 57.565 126.630 57.900 ;
        RECT 122.485 57.365 125.925 57.565 ;
        RECT 35.670 56.445 39.855 56.835 ;
        RECT 36.395 56.320 39.855 56.445 ;
        RECT 36.395 55.900 40.600 56.320 ;
        RECT 37.120 55.810 40.600 55.900 ;
        RECT 37.120 55.365 41.345 55.810 ;
        RECT 46.890 55.780 51.390 56.980 ;
        RECT 62.940 56.750 63.240 57.050 ;
        RECT 64.740 56.750 65.040 57.050 ;
        RECT 65.340 56.750 65.640 57.050 ;
        RECT 65.940 56.750 66.240 57.050 ;
        RECT 66.540 56.750 66.840 57.050 ;
        RECT 68.340 56.750 68.640 57.050 ;
        RECT 81.670 56.910 82.270 57.210 ;
        RECT 82.870 56.910 84.370 57.210 ;
        RECT 84.970 56.910 85.570 57.210 ;
        RECT 99.710 56.990 100.910 57.290 ;
        RECT 101.210 56.990 102.410 57.290 ;
        RECT 121.760 57.000 125.925 57.365 ;
        RECT 62.640 56.450 63.540 56.750 ;
        RECT 68.040 56.450 68.940 56.750 ;
        RECT 62.640 56.150 63.840 56.450 ;
        RECT 67.740 56.150 68.940 56.450 ;
        RECT 81.970 56.610 83.470 56.910 ;
        RECT 83.770 56.610 85.570 56.910 ;
        RECT 99.110 56.690 100.310 56.990 ;
        RECT 101.810 56.690 103.010 56.990 ;
        RECT 121.760 56.835 125.210 57.000 ;
        RECT 81.970 56.310 83.170 56.610 ;
        RECT 84.070 56.310 84.970 56.610 ;
        RECT 98.210 56.390 100.010 56.690 ;
        RECT 102.110 56.390 103.910 56.690 ;
        RECT 121.025 56.445 125.210 56.835 ;
        RECT 62.640 55.850 64.440 56.150 ;
        RECT 67.140 55.850 68.940 56.150 ;
        RECT 37.855 55.310 41.345 55.365 ;
        RECT 37.855 54.835 42.100 55.310 ;
        RECT 47.190 55.180 51.090 55.780 ;
        RECT 38.600 54.820 42.100 54.835 ;
        RECT 47.790 54.880 50.490 55.180 ;
        RECT 38.600 54.340 42.865 54.820 ;
        RECT 47.790 54.580 50.190 54.880 ;
        RECT 38.600 54.320 43.630 54.340 ;
        RECT 39.345 53.870 43.630 54.320 ;
        RECT 39.345 53.810 44.405 53.870 ;
        RECT 40.100 53.410 44.405 53.810 ;
        RECT 40.100 53.310 45.180 53.410 ;
        RECT 40.865 52.960 45.180 53.310 ;
        RECT 40.865 52.820 45.965 52.960 ;
        RECT 41.630 52.520 45.965 52.820 ;
        RECT 41.630 52.340 46.755 52.520 ;
        RECT 42.405 52.090 46.755 52.340 ;
        RECT 42.405 51.870 47.550 52.090 ;
        RECT 43.180 51.665 47.550 51.870 ;
        RECT 43.180 51.410 48.355 51.665 ;
        RECT 43.965 51.255 48.355 51.410 ;
        RECT 43.965 50.960 49.160 51.255 ;
        RECT 44.755 50.855 49.160 50.960 ;
        RECT 44.755 50.520 49.970 50.855 ;
        RECT 45.550 50.465 49.970 50.520 ;
        RECT 45.550 50.090 50.785 50.465 ;
        RECT 46.355 50.085 50.785 50.090 ;
        RECT 46.355 49.715 51.605 50.085 ;
        RECT 52.220 49.715 52.670 55.650 ;
        RECT 62.640 55.550 65.040 55.850 ;
        RECT 66.540 55.550 68.640 55.850 ;
        RECT 82.570 55.710 84.670 56.310 ;
        RECT 97.910 55.790 99.410 56.390 ;
        RECT 102.710 55.790 104.210 56.390 ;
        RECT 121.025 56.320 124.485 56.445 ;
        RECT 120.280 55.900 124.485 56.320 ;
        RECT 120.280 55.810 123.760 55.900 ;
        RECT 64.440 55.250 65.640 55.550 ;
        RECT 65.940 55.250 67.140 55.550 ;
        RECT 80.770 55.410 81.070 55.710 ;
        RECT 82.570 55.410 82.870 55.710 ;
        RECT 83.170 55.410 83.470 55.710 ;
        RECT 83.770 55.410 84.070 55.710 ;
        RECT 84.370 55.410 84.670 55.710 ;
        RECT 86.170 55.410 86.470 55.710 ;
        RECT 98.210 55.490 99.110 55.790 ;
        RECT 100.010 55.490 100.310 55.790 ;
        RECT 100.610 55.490 100.910 55.790 ;
        RECT 101.210 55.490 101.510 55.790 ;
        RECT 101.810 55.490 102.110 55.790 ;
        RECT 103.010 55.490 103.910 55.790 ;
        RECT 65.040 54.650 66.540 55.250 ;
        RECT 80.470 55.110 81.370 55.410 ;
        RECT 85.870 55.110 86.770 55.410 ;
        RECT 80.470 54.810 81.670 55.110 ;
        RECT 85.570 54.810 86.770 55.110 ;
        RECT 100.010 54.890 102.110 55.490 ;
        RECT 119.535 55.365 123.760 55.810 ;
        RECT 119.535 55.310 123.025 55.365 ;
        RECT 64.440 54.350 65.640 54.650 ;
        RECT 65.940 54.350 67.140 54.650 ;
        RECT 80.470 54.510 82.270 54.810 ;
        RECT 84.970 54.510 86.770 54.810 ;
        RECT 99.410 54.590 100.610 54.890 ;
        RECT 101.510 54.590 102.410 54.890 ;
        RECT 118.780 54.835 123.025 55.310 ;
        RECT 118.780 54.820 122.280 54.835 ;
        RECT 63.840 54.050 65.040 54.350 ;
        RECT 66.540 54.050 67.740 54.350 ;
        RECT 80.470 54.210 82.870 54.510 ;
        RECT 84.370 54.210 86.470 54.510 ;
        RECT 99.410 54.290 100.910 54.590 ;
        RECT 101.210 54.290 103.010 54.590 ;
        RECT 118.015 54.340 122.280 54.820 ;
        RECT 62.940 53.750 64.740 54.050 ;
        RECT 66.840 53.750 68.640 54.050 ;
        RECT 82.270 53.910 83.470 54.210 ;
        RECT 83.770 53.910 84.970 54.210 ;
        RECT 99.110 53.990 99.710 54.290 ;
        RECT 100.310 53.990 101.810 54.290 ;
        RECT 102.410 53.990 103.010 54.290 ;
        RECT 62.640 53.150 64.140 53.750 ;
        RECT 67.440 53.150 68.940 53.750 ;
        RECT 82.870 53.310 84.370 53.910 ;
        RECT 99.110 53.690 99.410 53.990 ;
        RECT 98.810 53.390 99.410 53.690 ;
        RECT 62.940 52.850 63.840 53.150 ;
        RECT 64.740 52.850 65.040 53.150 ;
        RECT 65.340 52.850 65.640 53.150 ;
        RECT 65.940 52.850 66.240 53.150 ;
        RECT 66.540 52.850 66.840 53.150 ;
        RECT 67.740 52.850 68.640 53.150 ;
        RECT 82.270 53.010 83.470 53.310 ;
        RECT 83.770 53.010 84.970 53.310 ;
        RECT 98.810 53.090 99.710 53.390 ;
        RECT 100.610 53.090 101.510 53.990 ;
        RECT 102.710 53.690 103.010 53.990 ;
        RECT 117.250 54.320 122.280 54.340 ;
        RECT 117.250 53.870 121.535 54.320 ;
        RECT 116.475 53.810 121.535 53.870 ;
        RECT 102.710 53.390 103.310 53.690 ;
        RECT 116.475 53.410 120.780 53.810 ;
        RECT 102.410 53.090 103.310 53.390 ;
        RECT 64.740 52.250 66.840 52.850 ;
        RECT 81.670 52.710 82.870 53.010 ;
        RECT 84.370 52.710 85.570 53.010 ;
        RECT 80.770 52.410 82.570 52.710 ;
        RECT 84.670 52.410 86.470 52.710 ;
        RECT 64.140 51.950 65.340 52.250 ;
        RECT 66.240 51.950 67.140 52.250 ;
        RECT 64.140 51.650 65.640 51.950 ;
        RECT 65.940 51.650 67.740 51.950 ;
        RECT 80.470 51.810 81.970 52.410 ;
        RECT 85.270 51.810 86.770 52.410 ;
        RECT 98.810 51.890 103.310 53.090 ;
        RECT 115.700 53.310 120.780 53.410 ;
        RECT 115.700 52.960 120.015 53.310 ;
        RECT 114.915 52.820 120.015 52.960 ;
        RECT 114.915 52.520 119.250 52.820 ;
        RECT 114.125 52.340 119.250 52.520 ;
        RECT 114.125 52.090 118.475 52.340 ;
        RECT 63.840 51.350 64.440 51.650 ;
        RECT 65.040 51.350 66.540 51.650 ;
        RECT 67.140 51.350 67.740 51.650 ;
        RECT 80.770 51.510 81.670 51.810 ;
        RECT 82.570 51.510 82.870 51.810 ;
        RECT 83.170 51.510 83.470 51.810 ;
        RECT 83.770 51.510 84.070 51.810 ;
        RECT 84.370 51.510 84.670 51.810 ;
        RECT 85.570 51.510 86.470 51.810 ;
        RECT 63.840 51.050 64.140 51.350 ;
        RECT 46.355 49.665 52.670 49.715 ;
        RECT 47.160 49.355 52.670 49.665 ;
        RECT 63.540 50.750 64.140 51.050 ;
        RECT 63.540 50.450 64.440 50.750 ;
        RECT 65.340 50.450 66.240 51.350 ;
        RECT 67.440 51.050 67.740 51.350 ;
        RECT 67.440 50.750 68.040 51.050 ;
        RECT 82.570 50.910 84.670 51.510 ;
        RECT 99.110 51.290 103.010 51.890 ;
        RECT 113.330 51.870 118.475 52.090 ;
        RECT 99.710 50.990 102.410 51.290 ;
        RECT 67.140 50.450 68.040 50.750 ;
        RECT 47.160 49.255 53.265 49.355 ;
        RECT 47.970 49.005 53.265 49.255 ;
        RECT 63.540 49.250 68.040 50.450 ;
        RECT 81.970 50.610 83.170 50.910 ;
        RECT 84.070 50.610 84.970 50.910 ;
        RECT 99.710 50.690 102.110 50.990 ;
        RECT 81.970 50.310 83.470 50.610 ;
        RECT 83.770 50.310 85.570 50.610 ;
        RECT 81.670 50.010 82.270 50.310 ;
        RECT 82.870 50.010 84.370 50.310 ;
        RECT 84.970 50.010 85.570 50.310 ;
        RECT 81.670 49.710 81.970 50.010 ;
        RECT 81.370 49.410 81.970 49.710 ;
        RECT 47.970 48.855 54.100 49.005 ;
        RECT 48.785 48.670 54.100 48.855 ;
        RECT 48.785 48.465 54.940 48.670 ;
        RECT 63.840 48.650 67.740 49.250 ;
        RECT 49.605 48.340 54.940 48.465 ;
        RECT 64.440 48.350 67.140 48.650 ;
        RECT 49.605 48.085 55.780 48.340 ;
        RECT 50.435 48.025 55.780 48.085 ;
        RECT 64.440 48.050 66.840 48.350 ;
        RECT 50.435 47.715 56.630 48.025 ;
        RECT 51.265 47.420 57.480 47.715 ;
        RECT 51.265 47.355 58.335 47.420 ;
        RECT 52.100 47.135 58.335 47.355 ;
        RECT 52.100 47.005 59.195 47.135 ;
        RECT 68.870 47.035 69.320 49.120 ;
        RECT 81.370 49.110 82.270 49.410 ;
        RECT 83.170 49.110 84.070 50.010 ;
        RECT 85.270 49.710 85.570 50.010 ;
        RECT 85.270 49.410 85.870 49.710 ;
        RECT 84.970 49.110 85.870 49.410 ;
        RECT 81.370 47.910 85.870 49.110 ;
        RECT 104.140 48.025 104.590 51.760 ;
        RECT 113.330 51.665 117.700 51.870 ;
        RECT 112.525 51.410 117.700 51.665 ;
        RECT 112.525 51.255 116.915 51.410 ;
        RECT 111.720 50.960 116.915 51.255 ;
        RECT 111.720 50.855 116.125 50.960 ;
        RECT 110.910 50.520 116.125 50.855 ;
        RECT 110.910 50.465 115.330 50.520 ;
        RECT 110.095 50.090 115.330 50.465 ;
        RECT 110.095 50.085 114.525 50.090 ;
        RECT 109.275 49.715 114.525 50.085 ;
        RECT 108.445 49.665 114.525 49.715 ;
        RECT 108.445 49.355 113.720 49.665 ;
        RECT 107.615 49.255 113.720 49.355 ;
        RECT 107.615 49.005 112.910 49.255 ;
        RECT 106.780 48.855 112.910 49.005 ;
        RECT 106.780 48.670 112.095 48.855 ;
        RECT 105.940 48.465 112.095 48.670 ;
        RECT 105.940 48.340 111.275 48.465 ;
        RECT 105.100 48.085 111.275 48.340 ;
        RECT 105.100 48.025 110.445 48.085 ;
        RECT 81.670 47.310 85.570 47.910 ;
        RECT 52.940 46.860 59.195 47.005 ;
        RECT 52.940 46.670 60.055 46.860 ;
        RECT 53.780 46.600 60.055 46.670 ;
        RECT 53.780 46.345 60.920 46.600 ;
        RECT 68.555 46.585 69.320 47.035 ;
        RECT 82.270 47.010 84.970 47.310 ;
        RECT 82.270 46.710 84.670 47.010 ;
        RECT 53.780 46.340 61.790 46.345 ;
        RECT 54.630 46.105 61.790 46.340 ;
        RECT 54.630 46.025 62.660 46.105 ;
        RECT 55.480 45.875 62.660 46.025 ;
        RECT 55.480 45.715 63.535 45.875 ;
        RECT 56.335 45.655 63.535 45.715 ;
        RECT 56.335 45.445 64.415 45.655 ;
        RECT 56.335 45.420 65.295 45.445 ;
        RECT 57.195 45.250 65.295 45.420 ;
        RECT 57.195 45.135 66.180 45.250 ;
        RECT 58.055 45.065 66.180 45.135 ;
        RECT 58.055 44.890 67.065 45.065 ;
        RECT 58.055 44.860 67.950 44.890 ;
        RECT 58.920 44.725 67.950 44.860 ;
        RECT 68.555 44.725 69.005 46.585 ;
        RECT 58.920 44.600 69.005 44.725 ;
        RECT 59.790 44.570 69.005 44.600 ;
        RECT 59.790 44.430 69.735 44.570 ;
        RECT 59.790 44.345 70.625 44.430 ;
        RECT 60.660 44.300 70.625 44.345 ;
        RECT 60.660 44.180 71.520 44.300 ;
        RECT 60.660 44.105 72.420 44.180 ;
        RECT 61.535 44.070 72.420 44.105 ;
        RECT 61.535 43.975 73.315 44.070 ;
        RECT 86.700 43.975 87.150 47.780 ;
        RECT 104.140 47.715 110.445 48.025 ;
        RECT 103.400 47.420 109.615 47.715 ;
        RECT 102.545 47.355 109.615 47.420 ;
        RECT 102.545 47.135 108.780 47.355 ;
        RECT 101.685 47.005 108.780 47.135 ;
        RECT 101.685 46.860 107.940 47.005 ;
        RECT 100.825 46.670 107.940 46.860 ;
        RECT 100.825 46.600 107.100 46.670 ;
        RECT 99.960 46.345 107.100 46.600 ;
        RECT 99.090 46.340 107.100 46.345 ;
        RECT 99.090 46.105 106.250 46.340 ;
        RECT 98.220 46.025 106.250 46.105 ;
        RECT 98.220 45.875 105.400 46.025 ;
        RECT 97.345 45.715 105.400 45.875 ;
        RECT 97.345 45.655 104.545 45.715 ;
        RECT 96.465 45.445 104.545 45.655 ;
        RECT 95.585 45.420 104.545 45.445 ;
        RECT 95.585 45.250 103.685 45.420 ;
        RECT 94.700 45.135 103.685 45.250 ;
        RECT 94.700 45.065 102.825 45.135 ;
        RECT 93.815 44.890 102.825 45.065 ;
        RECT 92.930 44.860 102.825 44.890 ;
        RECT 92.930 44.725 101.960 44.860 ;
        RECT 92.040 44.600 101.960 44.725 ;
        RECT 92.040 44.570 101.090 44.600 ;
        RECT 91.145 44.430 101.090 44.570 ;
        RECT 90.255 44.345 101.090 44.430 ;
        RECT 90.255 44.300 100.220 44.345 ;
        RECT 89.360 44.180 100.220 44.300 ;
        RECT 88.460 44.105 100.220 44.180 ;
        RECT 88.460 44.070 99.345 44.105 ;
        RECT 87.565 43.975 99.345 44.070 ;
        RECT 61.535 43.890 74.215 43.975 ;
        RECT 86.665 43.890 99.345 43.975 ;
        RECT 61.535 43.875 75.115 43.890 ;
        RECT 62.415 43.815 75.115 43.875 ;
        RECT 85.765 43.875 99.345 43.890 ;
        RECT 85.765 43.815 98.465 43.875 ;
        RECT 62.415 43.755 76.020 43.815 ;
        RECT 84.860 43.755 98.465 43.815 ;
        RECT 62.415 43.705 76.920 43.755 ;
        RECT 83.960 43.705 98.465 43.755 ;
        RECT 62.415 43.665 77.825 43.705 ;
        RECT 83.055 43.665 98.465 43.705 ;
        RECT 62.415 43.655 78.730 43.665 ;
        RECT 63.295 43.635 78.730 43.655 ;
        RECT 82.150 43.655 98.465 43.665 ;
        RECT 82.150 43.635 97.585 43.655 ;
        RECT 63.295 43.620 79.635 43.635 ;
        RECT 81.245 43.620 97.585 43.635 ;
        RECT 63.295 43.445 97.585 43.620 ;
        RECT 64.180 43.250 96.700 43.445 ;
        RECT 65.065 43.065 95.815 43.250 ;
        RECT 65.950 42.890 94.930 43.065 ;
        RECT 66.840 42.725 94.040 42.890 ;
        RECT 67.735 42.570 93.145 42.725 ;
        RECT 68.625 42.430 92.255 42.570 ;
        RECT 69.520 42.300 91.360 42.430 ;
        RECT 70.420 42.180 90.460 42.300 ;
        RECT 71.315 42.070 89.565 42.180 ;
        RECT 72.215 41.975 88.665 42.070 ;
        RECT 73.115 41.890 87.765 41.975 ;
        RECT 74.020 41.815 86.860 41.890 ;
        RECT 74.920 41.755 85.960 41.815 ;
        RECT 75.825 41.705 85.055 41.755 ;
        RECT 76.730 41.665 84.150 41.705 ;
        RECT 77.635 41.635 83.245 41.665 ;
        RECT 78.540 41.620 82.340 41.635 ;
        RECT 79.440 41.610 81.435 41.620 ;
      LAYER met3 ;
        RECT 85.810 223.665 86.230 224.265 ;
        RECT 88.570 223.665 88.990 224.265 ;
        RECT 91.330 223.665 91.750 224.265 ;
        RECT 91.720 221.360 92.300 221.370 ;
        RECT 90.300 219.400 90.800 220.000 ;
        RECT 61.410 218.030 62.100 218.730 ;
        RECT 91.560 217.050 92.560 221.360 ;
        RECT 3.120 216.050 92.560 217.050 ;
        RECT 3.240 216.040 4.340 216.050 ;
        RECT 59.930 215.430 60.780 215.750 ;
        RECT 60.050 215.420 60.700 215.430 ;
        RECT 52.150 214.660 52.750 215.210 ;
      LAYER met3 ;
        RECT 53.210 208.130 67.770 215.020 ;
        RECT 34.340 149.300 41.230 163.860 ;
        RECT 48.330 160.450 55.220 175.010 ;
        RECT 64.970 166.980 71.860 181.540 ;
        RECT 82.800 168.320 89.690 182.880 ;
        RECT 100.240 164.340 107.130 178.900 ;
        RECT 115.720 155.390 122.610 169.950 ;
      LAYER met3 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 68.170 149.600 91.570 152.200 ;
      LAYER met3 ;
        RECT 24.270 134.520 31.160 149.080 ;
      LAYER met3 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 60.370 134.000 99.370 144.400 ;
      LAYER met3 ;
        RECT 127.890 142.280 134.780 156.840 ;
        RECT 16.350 117.430 23.240 131.990 ;
      LAYER met3 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
      LAYER met3 ;
        RECT 133.000 126.170 139.890 140.730 ;
      LAYER met3 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 0.530 114.410 2.770 114.870 ;
        RECT 7.470 114.410 9.070 114.435 ;
        RECT 0.530 112.910 9.070 114.410 ;
        RECT 30.710 114.305 31.810 115.555 ;
        RECT 0.530 112.330 2.770 112.910 ;
        RECT 7.470 112.885 9.070 112.910 ;
      LAYER met3 ;
        RECT 19.000 99.550 25.890 114.110 ;
      LAYER met3 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
      LAYER met3 ;
        RECT 138.320 108.490 145.210 123.050 ;
      LAYER met3 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
      LAYER met3 ;
        RECT 21.620 82.460 28.510 97.020 ;
      LAYER met3 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
      LAYER met3 ;
        RECT 133.000 90.810 139.890 105.370 ;
      LAYER met3 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
      LAYER met3 ;
        RECT 31.690 65.360 38.580 79.920 ;
      LAYER met3 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
      LAYER met3 ;
        RECT 125.240 74.700 132.130 89.260 ;
        RECT 45.670 54.210 52.560 68.770 ;
        RECT 62.320 47.680 69.210 62.240 ;
        RECT 80.150 46.340 87.040 60.900 ;
        RECT 97.590 50.320 104.480 64.880 ;
        RECT 113.070 59.270 119.960 73.830 ;
      LAYER met4 ;
        RECT 30.670 223.050 30.970 224.760 ;
        RECT 33.430 223.050 33.730 224.760 ;
        RECT 36.190 223.050 36.490 224.760 ;
        RECT 38.950 223.050 39.250 224.760 ;
        RECT 41.710 223.050 42.010 224.760 ;
        RECT 44.470 223.050 44.770 224.760 ;
        RECT 47.230 223.050 47.530 224.760 ;
        RECT 49.990 223.050 50.290 224.760 ;
        RECT 52.750 223.050 53.050 224.760 ;
        RECT 55.510 223.050 55.810 224.760 ;
        RECT 58.270 223.050 58.570 224.760 ;
        RECT 61.030 223.050 61.330 224.760 ;
        RECT 63.790 223.050 64.090 224.760 ;
        RECT 66.550 223.050 66.850 224.760 ;
        RECT 69.310 223.050 69.610 224.760 ;
        RECT 72.070 223.050 72.370 224.760 ;
        RECT 74.830 223.050 75.130 224.760 ;
        RECT 77.590 223.050 77.890 224.760 ;
        RECT 80.350 223.050 80.650 224.760 ;
        RECT 83.110 223.050 83.410 224.760 ;
        RECT 85.870 224.095 86.170 224.760 ;
        RECT 88.630 224.095 88.930 224.760 ;
        RECT 91.390 224.095 91.690 224.760 ;
        RECT 85.855 223.685 86.185 224.095 ;
        RECT 88.615 223.685 88.945 224.095 ;
        RECT 91.375 223.685 91.705 224.095 ;
        RECT 1.000 222.050 83.410 223.050 ;
        RECT 94.150 222.110 94.450 224.760 ;
        RECT 1.000 220.760 2.500 222.050 ;
        RECT 52.375 215.190 52.725 222.050 ;
        RECT 60.490 218.650 61.490 222.050 ;
        RECT 90.410 221.810 94.450 222.110 ;
        RECT 90.410 220.000 90.710 221.810 ;
        RECT 90.300 219.400 90.800 220.000 ;
        RECT 60.490 218.140 62.030 218.650 ;
        RECT 61.490 218.110 62.030 218.140 ;
        RECT 90.410 217.570 90.710 219.400 ;
        RECT 60.170 217.270 90.710 217.570 ;
        RECT 60.170 215.755 60.470 217.270 ;
        RECT 59.975 215.425 60.735 215.755 ;
        RECT 52.195 214.685 52.725 215.190 ;
        RECT 52.195 214.680 52.705 214.685 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 68.170 149.600 91.570 152.200 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 60.370 134.000 99.370 144.400 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 0.575 112.325 1.000 114.875 ;
        RECT 2.500 112.325 2.690 114.875 ;
        RECT 6.500 114.110 31.920 115.610 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
  END
END tt_um_oscillating_bones
END LIBRARY

