* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VGND uo_out[0] uo_out[1] uo_out[3] VPWR
X0 a_13289_43697# uo_out[2].t2 VPWR.t69 VPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_16868_43697# a_17160_43997# a_17111_44089# VPWR.t77 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2 a_16596_43697# a_16868_43697# VGND.t59 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t73 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X4 VGND.t9 uo_out[0].t2 ring_0/skullfet_inverter_6.A VGND.t8 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X5 a_17360_43697# a_17160_43997# a_17509_43723# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6 VGND.t76 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND.t31 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t30 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X8 a_15221_43697# uo_out[1].t2 VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9 VPWR.t71 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X10 a_15179_44089# a_14664_43697# VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VGND.t37 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VGND.t36 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X12 ring_0/skullfet_inverter_6.A uo_out[0].t3 VPWR.t95 VPWR.t94 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X13 a_15577_43723# a_15357_43723# VGND.t40 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X14 VGND.t19 a_14664_43697# uo_out[2].t1 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR.t67 a_13289_43697# a_13296_43997# VPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 VGND.t80 a_15221_43697# a_15228_43997# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t51 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t50 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X18 a_13843_43723# a_13296_43997# a_13496_43697# VPWR.t103 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X19 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VPWR.t37 VPWR.t36 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X20 VGND.t79 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_8.A VGND.t78 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X21 a_16501_43697# a_16596_43697# VGND.t15 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X22 a_12637_43697# a_12732_43697# VPWR.t59 VPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X23 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t35 VGND.t34 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X24 VGND.t25 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t24 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X25 a_17289_43723# a_17153_43697# a_16868_43697# VPWR.t93 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 a_13224_43723# a_12732_43697# VGND.t48 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR.t21 a_14664_43697# uo_out[2].t0 VPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X29 VPWR.t99 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VPWR.t98 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X30 VGND.t63 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t62 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X31 a_17707_43723# a_17153_43697# a_17360_43697# VGND.t71 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X32 VGND.t61 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t60 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X33 a_15156_43723# a_14664_43697# VGND.t17 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X34 a_14936_43697# a_15228_43997# a_15179_44089# VPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X35 a_13289_43697# uo_out[2].t3 VGND.t53 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X36 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_7.A VPWR.t107 VPWR.t106 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X37 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VPWR.t31 VPWR.t30 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X38 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VPWR.t83 VPWR.t82 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X39 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_8.A VPWR.t53 VPWR.t52 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X40 VGND.t5 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X41 a_14664_43697# a_14936_43697# VGND.t23 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X42 a_15428_43697# a_15228_43997# a_15577_43723# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X43 VGND.t55 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X44 VGND.t77 a_13496_43697# a_13425_43723# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X45 a_13247_44089# a_12732_43697# VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X46 a_15221_43697# uo_out[1].t3 VGND.t7 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X47 a_16868_43697# a_17153_43697# a_17088_43723# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X48 a_13645_43723# a_13425_43723# VGND.t32 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X49 VPWR.t3 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VPWR.t2 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X50 VPWR.t35 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VPWR.t34 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X51 VGND.t69 a_15428_43697# a_15357_43723# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X52 VGND.t47 a_12732_43697# uo_out[3].t1 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 VGND.t11 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t10 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X54 VPWR.t75 a_17360_43697# a_17289_43723# VPWR.t74 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X55 a_14664_43697# a_14936_43697# VPWR.t29 VPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X56 VGND.t52 a_13289_43697# a_13296_43997# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X57 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VPWR.t81 VPWR.t80 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X58 VPWR.t43 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VPWR.t42 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X59 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X60 a_14569_43697# a_14664_43697# VGND.t16 VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X61 a_15604_44089# a_15357_43723# VPWR.t49 VPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X62 a_15357_43723# a_15221_43697# a_14936_43697# VPWR.t111 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X63 a_15428_43697# a_15221_43697# a_15604_44089# VPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X64 a_12732_43697# a_13004_43697# VGND.t21 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X65 VGND.t73 ring_0/skullfet_inverter_4.A uo_out[0].t1 VGND.t72 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X66 a_17289_43723# a_17160_43997# a_16868_43697# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X67 VPWR.t5 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X68 VPWR.t55 a_12732_43697# uo_out[3].t0 VPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X69 VGND.t67 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t66 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X70 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VPWR.t85 VPWR.t84 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X71 VPWR.t113 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VPWR.t112 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X72 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X73 a_17153_43697# uo_out[0].t4 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X74 a_17536_44089# a_17289_43723# VPWR.t1 VPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X75 a_15775_43723# a_15221_43697# a_15428_43697# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X76 a_17360_43697# a_17153_43697# a_17536_44089# VPWR.t92 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X77 a_17111_44089# a_16596_43697# VPWR.t17 VPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X78 a_13004_43697# a_13296_43997# a_13247_44089# VPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X79 VPWR.t61 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X80 a_12732_43697# a_13004_43697# VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X81 VGND.t42 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t41 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X82 VGND.t33 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X83 a_13496_43697# a_13296_43997# a_13645_43723# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X84 uo_out[0].t0 ring_0/skullfet_inverter_4.A VPWR.t97 VPWR.t96 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X85 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VPWR.t87 VPWR.t86 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X86 a_16501_43697# a_16596_43697# VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X87 a_14936_43697# a_15221_43697# a_15156_43723# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X88 VPWR.t91 a_17153_43697# a_17160_43997# VPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X89 VPWR.t89 a_15428_43697# a_15357_43723# VPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X90 VGND.t65 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t64 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X91 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VPWR.t51 VPWR.t50 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X92 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t82 VGND.t81 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X93 a_13425_43723# a_13296_43997# a_13004_43697# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X94 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VPWR.t47 VPWR.t46 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X95 a_12637_43697# a_12732_43697# VGND.t46 VGND.t45 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X96 a_13672_44089# a_13425_43723# VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X97 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X98 a_13425_43723# a_13289_43697# a_13004_43697# VPWR.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 a_13496_43697# a_13289_43697# a_13672_44089# VPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X100 VPWR.t101 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X101 a_15357_43723# a_15228_43997# a_14936_43697# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X102 VPWR.t41 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X103 VPWR.t33 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VPWR.t32 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X104 a_17153_43697# uo_out[0].t5 VGND.t22 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X105 a_13843_43723# a_13289_43697# a_13496_43697# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X106 a_17509_43723# a_17289_43723# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X107 VGND.t14 a_16596_43697# uo_out[1].t1 VGND.t13 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X108 a_13004_43697# a_13289_43697# a_13224_43723# VGND.t20 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X109 VGND.t57 a_17360_43697# a_17289_43723# VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X110 VGND.t49 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X111 VPWR.t109 a_15221_43697# a_15228_43997# VPWR.t108 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X112 VGND.t54 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X113 a_15775_43723# a_15228_43997# a_15428_43697# VPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X114 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X115 a_16596_43697# a_16868_43697# VPWR.t79 VPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X116 a_14569_43697# a_14664_43697# VPWR.t19 VPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X117 VGND.t39 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VGND.t38 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X118 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X119 a_17707_43723# a_17160_43997# a_17360_43697# VPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X120 VPWR.t13 a_16596_43697# uo_out[1].t0 VPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X121 VGND.t44 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_9.A VGND.t43 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X122 VPWR.t105 a_13496_43697# a_13425_43723# VPWR.t104 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X123 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VPWR.t63 VPWR.t62 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X124 VGND.t70 a_17153_43697# a_17160_43997# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X125 a_17088_43723# a_16596_43697# VGND.t12 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 uo_out[2].n2 uo_out[2].t0 313.104
R1 uo_out[2].n0 uo_out[2].t2 294.557
R2 uo_out[2].t1 uo_out[2].n2 265.769
R3 uo_out[2] uo_out[2].t1 262.318
R4 uo_out[2].n0 uo_out[2].t3 211.01
R5 uo_out[2].n1 uo_out[2].n0 152
R6 uo_out[2].n5 uo_out[2] 16.2155
R7 uo_out[2].n4 uo_out[2].n1 11.6311
R8 uo_out[2].n4 uo_out[2].n3 9.3005
R9 uo_out[2].n3 uo_out[2] 7.17626
R10 uo_out[2].n3 uo_out[2].n2 4.84898
R11 uo_out[2].n5 uo_out[2].n4 4.51042
R12 uo_out[2].n1 uo_out[2] 1.37896
R13 uo_out[2] uo_out[2].n5 0.0730806
R14 VPWR.n112 VPWR.t47 739.681
R15 VPWR.n114 VPWR.t35 739.681
R16 VPWR.n116 VPWR.t45 739.681
R17 VPWR.n150 VPWR.t37 739.681
R18 VPWR.n148 VPWR.t113 739.681
R19 VPWR.n84 VPWR.t87 739.681
R20 VPWR.n5 VPWR.t83 739.681
R21 VPWR.n85 VPWR.t33 739.681
R22 VPWR.n109 VPWR.t43 739.681
R23 VPWR.n122 VPWR.t3 739.681
R24 VPWR.n119 VPWR.t99 739.681
R25 VPWR.n153 VPWR.t31 739.681
R26 VPWR.n82 VPWR.t85 739.681
R27 VPWR.n80 VPWR.t53 739.681
R28 VPWR.n53 VPWR.t95 739.681
R29 VPWR.n30 VPWR.t97 739.681
R30 VPWR.n9 VPWR.t51 739.681
R31 VPWR.n6 VPWR.t63 739.681
R32 VPWR.n3 VPWR.t81 739.681
R33 VPWR.n56 VPWR.t11 739.681
R34 VPWR.n159 VPWR.t107 739.681
R35 VPWR.n112 VPWR.t46 707.852
R36 VPWR.n114 VPWR.t34 707.852
R37 VPWR.n116 VPWR.t44 707.852
R38 VPWR.n150 VPWR.t36 707.852
R39 VPWR.n148 VPWR.t112 707.852
R40 VPWR.n153 VPWR.t30 707.852
R41 VPWR.n84 VPWR.t86 707.852
R42 VPWR.n82 VPWR.t84 707.852
R43 VPWR.n80 VPWR.t52 707.852
R44 VPWR.n53 VPWR.t94 707.852
R45 VPWR.n30 VPWR.t96 707.852
R46 VPWR.n9 VPWR.t50 707.852
R47 VPWR.n6 VPWR.t62 707.852
R48 VPWR.n5 VPWR.t82 707.852
R49 VPWR.n3 VPWR.t80 707.852
R50 VPWR.n56 VPWR.t10 707.852
R51 VPWR.n159 VPWR.t106 707.852
R52 VPWR.n85 VPWR.t32 707.852
R53 VPWR.n109 VPWR.t42 707.852
R54 VPWR.n122 VPWR.t2 707.852
R55 VPWR.n119 VPWR.t98 707.852
R56 VPWR.n318 VPWR.t57 667.734
R57 VPWR.n286 VPWR.t23 667.734
R58 VPWR.n358 VPWR.t17 667.734
R59 VPWR.n333 VPWR.t71 666.677
R60 VPWR.n272 VPWR.t41 666.677
R61 VPWR.n238 VPWR.t5 666.677
R62 VPWR.t78 VPWR.t16 624.456
R63 VPWR.t22 VPWR.t28 624.456
R64 VPWR.t56 VPWR.t26 624.456
R65 VPWR.n336 VPWR.n335 604.394
R66 VPWR.n267 VPWR.n266 604.394
R67 VPWR.n376 VPWR.n375 604.394
R68 VPWR.t4 VPWR.t90 556.386
R69 VPWR.t14 VPWR.t12 556.386
R70 VPWR.t108 VPWR.t40 556.386
R71 VPWR.t20 VPWR.t18 556.386
R72 VPWR.t66 VPWR.t70 556.386
R73 VPWR.t54 VPWR.t58 556.386
R74 VPWR.n251 VPWR.t60 414.33
R75 VPWR.t100 VPWR.n342 414.33
R76 VPWR.t74 VPWR.t0 390.654
R77 VPWR.t48 VPWR.t88 390.654
R78 VPWR.t38 VPWR.t104 390.654
R79 VPWR.t16 VPWR.t77 337.384
R80 VPWR.t25 VPWR.t22 337.384
R81 VPWR.t102 VPWR.t56 337.384
R82 VPWR.n316 VPWR.n306 333.348
R83 VPWR.n288 VPWR.n258 333.348
R84 VPWR.n356 VPWR.n246 333.348
R85 VPWR.n302 VPWR.n301 320.976
R86 VPWR.n279 VPWR.n262 320.976
R87 VPWR.n243 VPWR.n242 320.976
R88 VPWR.t0 VPWR.t92 304.829
R89 VPWR.t110 VPWR.t48 304.829
R90 VPWR.t64 VPWR.t38 304.829
R91 VPWR.t60 VPWR.t14 287.072
R92 VPWR.t18 VPWR.t100 287.072
R93 VPWR.t58 VPWR.t72 287.072
R94 VPWR.t92 VPWR.t76 281.154
R95 VPWR.t93 VPWR.t74 281.154
R96 VPWR.t24 VPWR.t110 281.154
R97 VPWR.t88 VPWR.t111 281.154
R98 VPWR.t103 VPWR.t64 281.154
R99 VPWR.t104 VPWR.t65 281.154
R100 VPWR.n343 VPWR.n251 272.274
R101 VPWR.n343 VPWR 272.274
R102 VPWR.n342 VPWR.n341 272.274
R103 VPWR.n341 VPWR 272.274
R104 VPWR.t76 VPWR.t4 251.559
R105 VPWR.t40 VPWR.t24 251.559
R106 VPWR.t70 VPWR.t103 251.559
R107 VPWR.t90 VPWR.t6 248.599
R108 VPWR.t77 VPWR.t93 248.599
R109 VPWR.t12 VPWR.t78 248.599
R110 VPWR.t8 VPWR.t108 248.599
R111 VPWR.t111 VPWR.t25 248.599
R112 VPWR.t28 VPWR.t20 248.599
R113 VPWR.t68 VPWR.t66 248.599
R114 VPWR.t65 VPWR.t102 248.599
R115 VPWR.t26 VPWR.t54 248.599
R116 VPWR.n310 VPWR.n309 240.522
R117 VPWR.n294 VPWR.n255 240.522
R118 VPWR.n350 VPWR.n349 240.522
R119 VPWR.n341 VPWR.n340 213.119
R120 VPWR.n342 VPWR.n252 213.119
R121 VPWR.n344 VPWR.n343 213.119
R122 VPWR.n251 VPWR.n249 213.119
R123 VPWR.n301 VPWR.t39 113.98
R124 VPWR.n262 VPWR.t49 113.98
R125 VPWR.n242 VPWR.t1 113.98
R126 VPWR.t6 VPWR 91.745
R127 VPWR VPWR.t8 91.745
R128 VPWR VPWR.t68 91.745
R129 VPWR.n309 VPWR.t59 61.9872
R130 VPWR.n255 VPWR.t19 61.9872
R131 VPWR.n349 VPWR.t15 61.9872
R132 VPWR.n335 VPWR.t69 41.5552
R133 VPWR.n335 VPWR.t67 41.5552
R134 VPWR.n266 VPWR.t9 41.5552
R135 VPWR.n266 VPWR.t109 41.5552
R136 VPWR.n375 VPWR.t7 41.5552
R137 VPWR.n375 VPWR.t91 41.5552
R138 VPWR.n301 VPWR.t105 35.4605
R139 VPWR.n262 VPWR.t89 35.4605
R140 VPWR.n242 VPWR.t75 35.4605
R141 VPWR.n315 VPWR.n307 34.6358
R142 VPWR.n311 VPWR.n307 34.6358
R143 VPWR.n329 VPWR.n299 34.6358
R144 VPWR.n329 VPWR.n328 34.6358
R145 VPWR.n328 VPWR.n327 34.6358
R146 VPWR.n324 VPWR.n323 34.6358
R147 VPWR.n323 VPWR.n322 34.6358
R148 VPWR.n322 VPWR.n304 34.6358
R149 VPWR.n289 VPWR.n256 34.6358
R150 VPWR.n293 VPWR.n256 34.6358
R151 VPWR.n274 VPWR.n273 34.6358
R152 VPWR.n274 VPWR.n263 34.6358
R153 VPWR.n278 VPWR.n263 34.6358
R154 VPWR.n281 VPWR.n280 34.6358
R155 VPWR.n281 VPWR.n260 34.6358
R156 VPWR.n285 VPWR.n260 34.6358
R157 VPWR.n355 VPWR.n247 34.6358
R158 VPWR.n351 VPWR.n247 34.6358
R159 VPWR.n370 VPWR.n369 34.6358
R160 VPWR.n369 VPWR.n368 34.6358
R161 VPWR.n368 VPWR.n240 34.6358
R162 VPWR.n364 VPWR.n363 34.6358
R163 VPWR.n363 VPWR.n362 34.6358
R164 VPWR.n362 VPWR.n244 34.6358
R165 VPWR.n317 VPWR.n316 32.0005
R166 VPWR.n288 VPWR.n287 32.0005
R167 VPWR.n357 VPWR.n356 32.0005
R168 VPWR.n377 VPWR.n376 30.7593
R169 VPWR.n318 VPWR.n317 30.4946
R170 VPWR.n287 VPWR.n286 30.4946
R171 VPWR.n358 VPWR.n357 30.4946
R172 VPWR.n309 VPWR.t73 30.1692
R173 VPWR.n255 VPWR.t101 30.1692
R174 VPWR.n349 VPWR.t61 30.1692
R175 VPWR.n333 VPWR.n299 27.4829
R176 VPWR.n295 VPWR.n294 27.4829
R177 VPWR.n273 VPWR.n272 27.4829
R178 VPWR.n350 VPWR.n348 27.4829
R179 VPWR.n370 VPWR.n238 27.4829
R180 VPWR.n306 VPWR.t27 26.5955
R181 VPWR.n306 VPWR.t55 26.5955
R182 VPWR.n258 VPWR.t29 26.5955
R183 VPWR.n258 VPWR.t21 26.5955
R184 VPWR.n246 VPWR.t79 26.5955
R185 VPWR.n246 VPWR.t13 26.5955
R186 VPWR.n311 VPWR.n310 25.6005
R187 VPWR.n294 VPWR.n293 25.6005
R188 VPWR.n351 VPWR.n350 25.6005
R189 VPWR.n340 VPWR.n253 23.7181
R190 VPWR.n295 VPWR.n252 23.7181
R191 VPWR.n344 VPWR.n250 23.7181
R192 VPWR.n348 VPWR.n249 23.7181
R193 VPWR.n336 VPWR.n334 22.9652
R194 VPWR.n271 VPWR.n267 22.9652
R195 VPWR.n376 VPWR.n374 22.9652
R196 VPWR.n334 VPWR.n333 21.8358
R197 VPWR.n272 VPWR.n271 21.8358
R198 VPWR.n374 VPWR.n238 21.8358
R199 VPWR.n377 VPWR.n237 21.795
R200 VPWR.n336 VPWR.n253 21.4593
R201 VPWR.n267 VPWR.n250 21.4593
R202 VPWR.n327 VPWR.n302 18.4476
R203 VPWR.n279 VPWR.n278 18.4476
R204 VPWR.n243 VPWR.n240 18.4476
R205 VPWR.n324 VPWR.n302 16.1887
R206 VPWR.n280 VPWR.n279 16.1887
R207 VPWR.n364 VPWR.n243 16.1887
R208 VPWR.n318 VPWR.n304 15.0593
R209 VPWR.n286 VPWR.n285 15.0593
R210 VPWR.n358 VPWR.n244 15.0593
R211 VPWR.n154 VPWR.n153 13.377
R212 VPWR.n83 VPWR.n82 13.377
R213 VPWR.n81 VPWR.n80 13.377
R214 VPWR.n54 VPWR.n53 13.377
R215 VPWR.n31 VPWR.n30 13.377
R216 VPWR.n10 VPWR.n9 13.377
R217 VPWR.n7 VPWR.n6 13.377
R218 VPWR.n4 VPWR.n3 13.377
R219 VPWR.n57 VPWR.n56 13.377
R220 VPWR.n160 VPWR.n159 13.377
R221 VPWR VPWR.n112 13.3202
R222 VPWR.n115 VPWR.n114 13.3202
R223 VPWR VPWR.n116 13.3202
R224 VPWR VPWR.n150 13.3202
R225 VPWR.n149 VPWR.n148 13.3202
R226 VPWR VPWR.n84 13.3202
R227 VPWR VPWR.n5 13.3202
R228 VPWR.n86 VPWR.n85 13.3202
R229 VPWR.n110 VPWR.n109 13.3202
R230 VPWR.n123 VPWR.n122 13.3202
R231 VPWR.n120 VPWR.n119 13.3202
R232 VPWR.n340 VPWR.n252 12.8005
R233 VPWR.n344 VPWR.n249 12.8005
R234 VPWR.n113 VPWR 9.7375
R235 VPWR.n117 VPWR 9.39357
R236 VPWR.n376 VPWR.n0 9.3005
R237 VPWR.n374 VPWR.n373 9.3005
R238 VPWR.n372 VPWR.n238 9.3005
R239 VPWR.n371 VPWR.n370 9.3005
R240 VPWR.n369 VPWR.n239 9.3005
R241 VPWR.n368 VPWR.n367 9.3005
R242 VPWR.n366 VPWR.n240 9.3005
R243 VPWR.n365 VPWR.n364 9.3005
R244 VPWR.n363 VPWR.n241 9.3005
R245 VPWR.n362 VPWR.n361 9.3005
R246 VPWR.n360 VPWR.n244 9.3005
R247 VPWR.n359 VPWR.n358 9.3005
R248 VPWR.n357 VPWR.n245 9.3005
R249 VPWR.n355 VPWR.n354 9.3005
R250 VPWR.n353 VPWR.n247 9.3005
R251 VPWR.n352 VPWR.n351 9.3005
R252 VPWR.n350 VPWR.n248 9.3005
R253 VPWR.n348 VPWR.n347 9.3005
R254 VPWR.n346 VPWR.n249 9.3005
R255 VPWR.n345 VPWR.n344 9.3005
R256 VPWR.n268 VPWR.n250 9.3005
R257 VPWR.n269 VPWR.n267 9.3005
R258 VPWR.n271 VPWR.n270 9.3005
R259 VPWR.n272 VPWR.n265 9.3005
R260 VPWR.n273 VPWR.n264 9.3005
R261 VPWR.n275 VPWR.n274 9.3005
R262 VPWR.n276 VPWR.n263 9.3005
R263 VPWR.n278 VPWR.n277 9.3005
R264 VPWR.n280 VPWR.n261 9.3005
R265 VPWR.n282 VPWR.n281 9.3005
R266 VPWR.n283 VPWR.n260 9.3005
R267 VPWR.n285 VPWR.n284 9.3005
R268 VPWR.n286 VPWR.n259 9.3005
R269 VPWR.n287 VPWR.n257 9.3005
R270 VPWR.n290 VPWR.n289 9.3005
R271 VPWR.n291 VPWR.n256 9.3005
R272 VPWR.n293 VPWR.n292 9.3005
R273 VPWR.n294 VPWR.n254 9.3005
R274 VPWR.n296 VPWR.n295 9.3005
R275 VPWR.n297 VPWR.n252 9.3005
R276 VPWR.n340 VPWR.n339 9.3005
R277 VPWR.n338 VPWR.n253 9.3005
R278 VPWR.n337 VPWR.n336 9.3005
R279 VPWR.n334 VPWR.n298 9.3005
R280 VPWR.n333 VPWR.n332 9.3005
R281 VPWR.n331 VPWR.n299 9.3005
R282 VPWR.n330 VPWR.n329 9.3005
R283 VPWR.n328 VPWR.n300 9.3005
R284 VPWR.n327 VPWR.n326 9.3005
R285 VPWR.n325 VPWR.n324 9.3005
R286 VPWR.n323 VPWR.n303 9.3005
R287 VPWR.n322 VPWR.n321 9.3005
R288 VPWR.n320 VPWR.n304 9.3005
R289 VPWR.n319 VPWR.n318 9.3005
R290 VPWR.n317 VPWR.n305 9.3005
R291 VPWR.n315 VPWR.n314 9.3005
R292 VPWR.n313 VPWR.n307 9.3005
R293 VPWR.n312 VPWR.n311 9.3005
R294 VPWR.n155 VPWR.n154 8.51977
R295 VPWR.n232 VPWR 8.13646
R296 VPWR.n121 VPWR.n118 7.53241
R297 VPWR.n157 VPWR.n83 7.53109
R298 VPWR.n158 VPWR.n81 7.45619
R299 VPWR.n310 VPWR.n308 7.4049
R300 VPWR.n151 VPWR 7.19357
R301 VPWR.n161 VPWR.n160 6.79323
R302 VPWR.n233 VPWR.n4 6.76538
R303 VPWR.n156 VPWR 6.40107
R304 VPWR.n121 VPWR.n120 6.34337
R305 VPWR.n124 VPWR.n123 6.19552
R306 VPWR.n117 VPWR.n115 6.1805
R307 VPWR.n231 VPWR.n7 6.08268
R308 VPWR.n118 VPWR.n113 6.07746
R309 VPWR.n58 VPWR.n57 6.01772
R310 VPWR.n229 VPWR.n10 6.01019
R311 VPWR.n32 VPWR.n31 5.71852
R312 VPWR.n55 VPWR.n54 5.65925
R313 VPWR.n111 VPWR.n110 5.44488
R314 VPWR.n87 VPWR.n86 5.3655
R315 VPWR.n151 VPWR.n149 5.233
R316 VPWR.n231 VPWR.n230 4.17361
R317 VPWR.n155 VPWR.n152 4.09662
R318 VPWR.n237 VPWR 3.1965
R319 VPWR.n186 VPWR.n185 3.07281
R320 VPWR.n316 VPWR.n315 2.63579
R321 VPWR.n289 VPWR.n288 2.63579
R322 VPWR.n356 VPWR.n355 2.63579
R323 VPWR.n237 VPWR.n236 1.96192
R324 VPWR.n118 VPWR.n117 1.25038
R325 VPWR.n152 VPWR.n147 1.04638
R326 VPWR.n156 VPWR.n155 0.926193
R327 VPWR.n124 VPWR.n121 0.897709
R328 VPWR.n157 VPWR.n156 0.877511
R329 VPWR.n224 VPWR.n223 0.861295
R330 VPWR.n232 VPWR.n231 0.838747
R331 VPWR.n233 VPWR.n232 0.810795
R332 VPWR.n113 VPWR.n2 0.786394
R333 VPWR.n162 VPWR.n158 0.69817
R334 VPWR.n125 VPWR.n124 0.574375
R335 VPWR.n158 VPWR.n157 0.53698
R336 VPWR.n225 VPWR.n224 0.507602
R337 VPWR.n185 VPWR.n184 0.491158
R338 VPWR.n152 VPWR.n151 0.456575
R339 VPWR.n226 VPWR.n225 0.391496
R340 VPWR.n187 VPWR.n186 0.380996
R341 VPWR.n235 VPWR.n234 0.341219
R342 VPWR.n226 VPWR.n8 0.325974
R343 VPWR.n125 VPWR.n111 0.323617
R344 VPWR.n230 VPWR.n8 0.320751
R345 VPWR.n188 VPWR.n187 0.263105
R346 VPWR.n189 VPWR.n188 0.23221
R347 VPWR.n228 VPWR.n8 0.198913
R348 VPWR.n227 VPWR.n226 0.195812
R349 VPWR.n190 VPWR.n189 0.193814
R350 VPWR.n225 VPWR.n11 0.192808
R351 VPWR.n224 VPWR.n12 0.189894
R352 VPWR.n235 VPWR.n2 0.188146
R353 VPWR.n191 VPWR.n190 0.183989
R354 VPWR.n163 VPWR.n162 0.169675
R355 VPWR.n184 VPWR.n183 0.168706
R356 VPWR.n186 VPWR.n52 0.162658
R357 VPWR.n192 VPWR.n191 0.157627
R358 VPWR.n308 VPWR 0.156264
R359 VPWR.n14 VPWR.n13 0.154418
R360 VPWR.n161 VPWR.n79 0.154418
R361 VPWR.n208 VPWR.n28 0.153485
R362 VPWR.n193 VPWR.n192 0.148565
R363 VPWR.n89 VPWR.n88 0.147626
R364 VPWR.n312 VPWR.n308 0.144904
R365 VPWR.n187 VPWR.n51 0.143882
R366 VPWR.n188 VPWR.n50 0.142412
R367 VPWR.n190 VPWR.n48 0.140206
R368 VPWR.n189 VPWR.n49 0.140035
R369 VPWR.n192 VPWR.n46 0.139637
R370 VPWR.n191 VPWR.n47 0.139471
R371 VPWR.n127 VPWR.n107 0.137548
R372 VPWR.n194 VPWR.n44 0.137405
R373 VPWR.n193 VPWR.n45 0.137265
R374 VPWR.n129 VPWR.n105 0.136933
R375 VPWR.n195 VPWR.n43 0.136661
R376 VPWR.n126 VPWR.n108 0.136661
R377 VPWR.n221 VPWR.n15 0.136529
R378 VPWR.n164 VPWR.n78 0.136529
R379 VPWR.n128 VPWR.n106 0.136042
R380 VPWR.n196 VPWR.n42 0.135917
R381 VPWR.n194 VPWR.n193 0.135794
R382 VPWR.n182 VPWR.n60 0.135785
R383 VPWR.n144 VPWR.n90 0.135774
R384 VPWR.n133 VPWR.n101 0.135656
R385 VPWR.n222 VPWR.n14 0.13561
R386 VPWR.n163 VPWR.n79 0.13561
R387 VPWR.n132 VPWR.n102 0.135531
R388 VPWR.n130 VPWR.n104 0.135409
R389 VPWR.n140 VPWR.n94 0.135368
R390 VPWR.n219 VPWR.n17 0.135321
R391 VPWR.n166 VPWR.n76 0.135321
R392 VPWR.n198 VPWR.n40 0.135289
R393 VPWR.n138 VPWR.n96 0.13524
R394 VPWR.n135 VPWR.n99 0.134994
R395 VPWR.n145 VPWR.n89 0.134918
R396 VPWR.n142 VPWR.n92 0.134667
R397 VPWR.n197 VPWR.n41 0.134429
R398 VPWR.n136 VPWR.n98 0.134203
R399 VPWR.n201 VPWR.n37 0.133884
R400 VPWR.n200 VPWR.n38 0.133884
R401 VPWR.n131 VPWR.n103 0.133884
R402 VPWR.n199 VPWR.n39 0.133783
R403 VPWR.n209 VPWR.n27 0.133617
R404 VPWR.n176 VPWR.n66 0.133617
R405 VPWR.n220 VPWR.n16 0.133536
R406 VPWR.n165 VPWR.n77 0.133536
R407 VPWR.n217 VPWR.n19 0.133312
R408 VPWR.n204 VPWR.n34 0.133312
R409 VPWR.n181 VPWR.n61 0.133312
R410 VPWR.n168 VPWR.n74 0.133312
R411 VPWR.n215 VPWR.n21 0.133205
R412 VPWR.n171 VPWR.n71 0.133101
R413 VPWR.n143 VPWR.n91 0.133
R414 VPWR.n211 VPWR.n25 0.132901
R415 VPWR.n174 VPWR.n68 0.132901
R416 VPWR.n141 VPWR.n93 0.132901
R417 VPWR.n206 VPWR.n32 0.13262
R418 VPWR.n179 VPWR.n63 0.13262
R419 VPWR.n137 VPWR.n97 0.13262
R420 VPWR.n203 VPWR.n35 0.132444
R421 VPWR.n134 VPWR.n100 0.132444
R422 VPWR.n202 VPWR.n36 0.13236
R423 VPWR.n216 VPWR.n20 0.132349
R424 VPWR.n169 VPWR.n73 0.132349
R425 VPWR.n213 VPWR.n23 0.132167
R426 VPWR.n172 VPWR.n70 0.132167
R427 VPWR.n139 VPWR.n95 0.13191
R428 VPWR.n178 VPWR.n64 0.131829
R429 VPWR.n108 VPWR.n107 0.131701
R430 VPWR.n218 VPWR.n18 0.131576
R431 VPWR.n167 VPWR.n75 0.131576
R432 VPWR.n170 VPWR.n72 0.131412
R433 VPWR.n214 VPWR.n22 0.131333
R434 VPWR.n212 VPWR.n24 0.131257
R435 VPWR.n173 VPWR.n69 0.131257
R436 VPWR.n205 VPWR.n33 0.130901
R437 VPWR.n180 VPWR.n62 0.130901
R438 VPWR.n147 VPWR.n146 0.130756
R439 VPWR.n177 VPWR.n65 0.130247
R440 VPWR.n107 VPWR.n106 0.130144
R441 VPWR.n195 VPWR.n194 0.130052
R442 VPWR.n210 VPWR.n26 0.129506
R443 VPWR.n175 VPWR.n67 0.129506
R444 VPWR.n183 VPWR.n59 0.12922
R445 VPWR.n222 VPWR.n221 0.124945
R446 VPWR.n164 VPWR.n163 0.124945
R447 VPWR.n196 VPWR.n195 0.12426
R448 VPWR.n221 VPWR.n220 0.122959
R449 VPWR.n165 VPWR.n164 0.122959
R450 VPWR.n106 VPWR.n105 0.122756
R451 VPWR.n105 VPWR.n104 0.122197
R452 VPWR.n208 VPWR.n207 0.121074
R453 VPWR.n373 VPWR.n0 0.120292
R454 VPWR.n373 VPWR.n372 0.120292
R455 VPWR.n372 VPWR.n371 0.120292
R456 VPWR.n371 VPWR.n239 0.120292
R457 VPWR.n367 VPWR.n239 0.120292
R458 VPWR.n367 VPWR.n366 0.120292
R459 VPWR.n366 VPWR.n365 0.120292
R460 VPWR.n365 VPWR.n241 0.120292
R461 VPWR.n361 VPWR.n241 0.120292
R462 VPWR.n361 VPWR.n360 0.120292
R463 VPWR.n360 VPWR.n359 0.120292
R464 VPWR.n359 VPWR.n245 0.120292
R465 VPWR.n354 VPWR.n245 0.120292
R466 VPWR.n354 VPWR.n353 0.120292
R467 VPWR.n353 VPWR.n352 0.120292
R468 VPWR.n352 VPWR.n248 0.120292
R469 VPWR.n347 VPWR.n248 0.120292
R470 VPWR.n270 VPWR.n269 0.120292
R471 VPWR.n270 VPWR.n265 0.120292
R472 VPWR.n265 VPWR.n264 0.120292
R473 VPWR.n275 VPWR.n264 0.120292
R474 VPWR.n276 VPWR.n275 0.120292
R475 VPWR.n277 VPWR.n276 0.120292
R476 VPWR.n277 VPWR.n261 0.120292
R477 VPWR.n282 VPWR.n261 0.120292
R478 VPWR.n283 VPWR.n282 0.120292
R479 VPWR.n284 VPWR.n283 0.120292
R480 VPWR.n284 VPWR.n259 0.120292
R481 VPWR.n259 VPWR.n257 0.120292
R482 VPWR.n290 VPWR.n257 0.120292
R483 VPWR.n291 VPWR.n290 0.120292
R484 VPWR.n292 VPWR.n291 0.120292
R485 VPWR.n292 VPWR.n254 0.120292
R486 VPWR.n296 VPWR.n254 0.120292
R487 VPWR.n337 VPWR.n298 0.120292
R488 VPWR.n332 VPWR.n298 0.120292
R489 VPWR.n332 VPWR.n331 0.120292
R490 VPWR.n331 VPWR.n330 0.120292
R491 VPWR.n330 VPWR.n300 0.120292
R492 VPWR.n326 VPWR.n300 0.120292
R493 VPWR.n326 VPWR.n325 0.120292
R494 VPWR.n325 VPWR.n303 0.120292
R495 VPWR.n321 VPWR.n303 0.120292
R496 VPWR.n321 VPWR.n320 0.120292
R497 VPWR.n320 VPWR.n319 0.120292
R498 VPWR.n319 VPWR.n305 0.120292
R499 VPWR.n314 VPWR.n305 0.120292
R500 VPWR.n314 VPWR.n313 0.120292
R501 VPWR.n313 VPWR.n312 0.120292
R502 VPWR.n220 VPWR.n219 0.12023
R503 VPWR.n166 VPWR.n165 0.12023
R504 VPWR.n219 VPWR.n218 0.119565
R505 VPWR.n167 VPWR.n166 0.119565
R506 VPWR.n228 VPWR.n227 0.118556
R507 VPWR.n147 VPWR.n87 0.118474
R508 VPWR.n104 VPWR.n103 0.117381
R509 VPWR.n197 VPWR.n196 0.117018
R510 VPWR.n198 VPWR.n197 0.116571
R511 VPWR.n218 VPWR.n217 0.115278
R512 VPWR.n168 VPWR.n167 0.115278
R513 VPWR.n227 VPWR.n11 0.114758
R514 VPWR.n90 VPWR.n89 0.114696
R515 VPWR.n207 VPWR.n29 0.114511
R516 VPWR.n217 VPWR.n216 0.114352
R517 VPWR.n169 VPWR.n168 0.114352
R518 VPWR.n102 VPWR.n101 0.114094
R519 VPWR.n216 VPWR.n215 0.113756
R520 VPWR.n170 VPWR.n169 0.113235
R521 VPWR.n92 VPWR.n91 0.113192
R522 VPWR.n101 VPWR.n100 0.113154
R523 VPWR.n91 VPWR.n90 0.112678
R524 VPWR.n94 VPWR.n93 0.112433
R525 VPWR.n209 VPWR.n208 0.112207
R526 VPWR.n199 VPWR.n198 0.111422
R527 VPWR.n215 VPWR.n214 0.111333
R528 VPWR.n98 VPWR.n97 0.111285
R529 VPWR.n214 VPWR.n213 0.111081
R530 VPWR.n172 VPWR.n171 0.111081
R531 VPWR.n12 VPWR.n11 0.111077
R532 VPWR.n171 VPWR.n170 0.110429
R533 VPWR.n96 VPWR.n95 0.110229
R534 VPWR.n173 VPWR.n172 0.11011
R535 VPWR.n93 VPWR.n92 0.109923
R536 VPWR.n103 VPWR.n102 0.10979
R537 VPWR.n201 VPWR.n200 0.109555
R538 VPWR.n183 VPWR.n182 0.108951
R539 VPWR.n211 VPWR.n210 0.108673
R540 VPWR.n175 VPWR.n174 0.108673
R541 VPWR.n213 VPWR.n212 0.108622
R542 VPWR.n99 VPWR.n98 0.108359
R543 VPWR.n100 VPWR.n99 0.108286
R544 VPWR.n95 VPWR.n94 0.10823
R545 VPWR.n200 VPWR.n199 0.107819
R546 VPWR.n97 VPWR.n96 0.107643
R547 VPWR.n236 VPWR.n235 0.107643
R548 VPWR.n212 VPWR.n211 0.107267
R549 VPWR.n174 VPWR.n173 0.107267
R550 VPWR.n177 VPWR.n176 0.107106
R551 VPWR.n13 VPWR.n12 0.106561
R552 VPWR.n202 VPWR.n201 0.105203
R553 VPWR.n203 VPWR.n202 0.105131
R554 VPWR.n182 VPWR.n181 0.104693
R555 VPWR.n205 VPWR.n204 0.104583
R556 VPWR.n181 VPWR.n180 0.104583
R557 VPWR.n204 VPWR.n203 0.104127
R558 VPWR.n206 VPWR.n205 0.103965
R559 VPWR.n180 VPWR.n179 0.103965
R560 VPWR.n207 VPWR.n206 0.103813
R561 VPWR.n179 VPWR.n178 0.103813
R562 VPWR.n178 VPWR.n177 0.103788
R563 VPWR.n210 VPWR.n209 0.103439
R564 VPWR.n176 VPWR.n175 0.103439
R565 VPWR.n223 VPWR.n222 0.100519
R566 VPWR VPWR.n0 0.0981562
R567 VPWR.n269 VPWR 0.0981562
R568 VPWR VPWR.n337 0.0981562
R569 VPWR.n15 VPWR.n14 0.0979265
R570 VPWR.n79 VPWR.n78 0.0979265
R571 VPWR.n16 VPWR.n15 0.0960882
R572 VPWR.n78 VPWR.n77 0.0960882
R573 VPWR.n17 VPWR.n16 0.0915714
R574 VPWR.n77 VPWR.n76 0.0915714
R575 VPWR.n18 VPWR.n17 0.088
R576 VPWR.n76 VPWR.n75 0.088
R577 VPWR.n19 VPWR.n18 0.0855694
R578 VPWR.n75 VPWR.n74 0.0855694
R579 VPWR.n146 VPWR.n88 0.0849982
R580 VPWR.n223 VPWR.n13 0.0844552
R581 VPWR.n230 VPWR.n229 0.0832089
R582 VPWR.n20 VPWR.n19 0.0820972
R583 VPWR.n74 VPWR.n73 0.0820972
R584 VPWR.n21 VPWR.n20 0.0792671
R585 VPWR.n73 VPWR.n72 0.0792671
R586 VPWR.n22 VPWR.n21 0.0775548
R587 VPWR.n72 VPWR.n71 0.0765135
R588 VPWR.n146 VPWR.n145 0.0741301
R589 VPWR.n71 VPWR.n70 0.0731351
R590 VPWR.n145 VPWR.n144 0.0724178
R591 VPWR.n23 VPWR.n22 0.0721667
R592 VPWR.n24 VPWR.n23 0.0705
R593 VPWR.n70 VPWR.n69 0.0705
R594 VPWR.n144 VPWR.n143 0.0688333
R595 VPWR.n25 VPWR.n24 0.0679342
R596 VPWR.n69 VPWR.n68 0.0679342
R597 VPWR.n29 VPWR.n28 0.0676642
R598 VPWR.n143 VPWR.n142 0.0655
R599 VPWR.n26 VPWR.n25 0.0646447
R600 VPWR.n68 VPWR.n67 0.0646447
R601 VPWR.n142 VPWR.n141 0.0646447
R602 VPWR.n27 VPWR.n26 0.063
R603 VPWR.n67 VPWR.n66 0.063
R604 VPWR.n347 VPWR 0.0603958
R605 VPWR VPWR.n346 0.0603958
R606 VPWR VPWR.n345 0.0603958
R607 VPWR.n268 VPWR 0.0603958
R608 VPWR VPWR.n296 0.0603958
R609 VPWR.n297 VPWR 0.0603958
R610 VPWR.n339 VPWR 0.0603958
R611 VPWR VPWR.n338 0.0603958
R612 VPWR.n141 VPWR.n140 0.0597105
R613 VPWR.n28 VPWR.n27 0.0589416
R614 VPWR.n66 VPWR.n65 0.0589416
R615 VPWR.n140 VPWR.n139 0.0581923
R616 VPWR.n65 VPWR.n64 0.057462
R617 VPWR.n154 VPWR 0.0573182
R618 VPWR.n83 VPWR 0.0573182
R619 VPWR.n81 VPWR 0.0573182
R620 VPWR.n54 VPWR 0.0573182
R621 VPWR.n31 VPWR 0.0573182
R622 VPWR.n10 VPWR 0.0573182
R623 VPWR.n7 VPWR 0.0573182
R624 VPWR.n4 VPWR 0.0573182
R625 VPWR.n57 VPWR 0.0573182
R626 VPWR.n160 VPWR 0.0573182
R627 VPWR.n139 VPWR.n138 0.0556948
R628 VPWR.n64 VPWR.n63 0.0542975
R629 VPWR.n33 VPWR.n32 0.0527152
R630 VPWR.n63 VPWR.n62 0.0527152
R631 VPWR.n138 VPWR.n137 0.0527152
R632 VPWR.n115 VPWR 0.0505
R633 VPWR.n149 VPWR 0.0505
R634 VPWR.n86 VPWR 0.0505
R635 VPWR.n110 VPWR 0.0505
R636 VPWR.n123 VPWR 0.0505
R637 VPWR.n120 VPWR 0.0505
R638 VPWR.n137 VPWR.n136 0.0495506
R639 VPWR.n34 VPWR.n33 0.0483395
R640 VPWR.n62 VPWR.n61 0.0483395
R641 VPWR.n136 VPWR.n135 0.0479684
R642 VPWR.n35 VPWR.n34 0.047375
R643 VPWR.n61 VPWR.n60 0.047375
R644 VPWR.n32 VPWR.n29 0.0472033
R645 VPWR.n60 VPWR.n59 0.0463861
R646 VPWR.n36 VPWR.n35 0.0452531
R647 VPWR.n135 VPWR.n134 0.0452531
R648 VPWR.n134 VPWR.n133 0.0426875
R649 VPWR.n37 VPWR.n36 0.0416585
R650 VPWR.n59 VPWR.n58 0.0406786
R651 VPWR.n88 VPWR.n87 0.039507
R652 VPWR.n133 VPWR.n132 0.0390802
R653 VPWR.n38 VPWR.n37 0.0386098
R654 VPWR.n39 VPWR.n38 0.0386098
R655 VPWR.n132 VPWR.n131 0.0386098
R656 VPWR.n346 VPWR 0.0382604
R657 VPWR.n345 VPWR 0.0382604
R658 VPWR VPWR.n297 0.0382604
R659 VPWR.n339 VPWR 0.0382604
R660 VPWR.n131 VPWR.n130 0.035561
R661 VPWR.n40 VPWR.n39 0.0351386
R662 VPWR.n126 VPWR.n125 0.0350681
R663 VPWR.n130 VPWR.n129 0.0325122
R664 VPWR.n41 VPWR.n40 0.0321265
R665 VPWR.n129 VPWR.n128 0.0306205
R666 VPWR.n42 VPWR.n41 0.0302619
R667 VPWR.n128 VPWR.n127 0.0276084
R668 VPWR.n43 VPWR.n42 0.0272857
R669 VPWR.n44 VPWR.n43 0.0257976
R670 VPWR.n127 VPWR.n126 0.0257976
R671 VPWR.n55 VPWR.n52 0.0244583
R672 VPWR.n45 VPWR.n44 0.0243095
R673 VPWR.n236 VPWR.n1 0.0243095
R674 VPWR.n185 VPWR.n55 0.0239375
R675 VPWR.n184 VPWR.n58 0.0227865
R676 VPWR VPWR.n268 0.0226354
R677 VPWR.n338 VPWR 0.0226354
R678 VPWR VPWR.n377 0.0224072
R679 VPWR.n2 VPWR.n1 0.0214028
R680 VPWR.n46 VPWR.n45 0.0210882
R681 VPWR.n47 VPWR.n46 0.0198452
R682 VPWR.n48 VPWR.n47 0.0166765
R683 VPWR.n49 VPWR.n48 0.0152059
R684 VPWR.n234 VPWR.n233 0.01479
R685 VPWR.n111 VPWR.n108 0.0131488
R686 VPWR.n234 VPWR.n1 0.0124293
R687 VPWR.n50 VPWR.n49 0.0121279
R688 VPWR.n51 VPWR.n50 0.0107941
R689 VPWR.n162 VPWR.n161 0.0104434
R690 VPWR.n52 VPWR.n51 0.00785294
R691 VPWR.n229 VPWR.n228 0.00590163
R692 VGND.n441 VGND.n62 171881
R693 VGND.n459 VGND.n458 156689
R694 VGND.n65 VGND.t24 151322
R695 VGND.n438 VGND.n75 130569
R696 VGND.n485 VGND.n484 130542
R697 VGND.n118 VGND.n72 49690.4
R698 VGND.n126 VGND.n3 48636.9
R699 VGND.n444 VGND.n75 45450.3
R700 VGND.n486 VGND.n485 44132.5
R701 VGND.n438 VGND.n437 44106
R702 VGND.n439 VGND.n77 43377.2
R703 VGND.n437 VGND.t10 31560.8
R704 VGND.n487 VGND.n486 30151.8
R705 VGND.n437 VGND.n77 29891.4
R706 VGND.n486 VGND.n1 29891.4
R707 VGND.n306 VGND.t58 18687.3
R708 VGND.n444 VGND.n62 16600.2
R709 VGND.n136 VGND.n131 16072.7
R710 VGND.n76 VGND.n61 14081.5
R711 VGND.n309 VGND.n118 13406.4
R712 VGND.n306 VGND.n305 13301.5
R713 VGND.n121 VGND.n120 12272.6
R714 VGND.n144 VGND.n121 12077.4
R715 VGND.n445 VGND.n444 11373.6
R716 VGND.n439 VGND.n438 10649.3
R717 VGND.n485 VGND.n3 10649.2
R718 VGND.n444 VGND.n72 8289.38
R719 VGND.n123 VGND.n121 6135.59
R720 VGND.n440 VGND.n439 6127.89
R721 VGND.n306 VGND 5326.64
R722 VGND.n309 VGND.n119 4245.54
R723 VGND.t60 VGND.n135 4169.04
R724 VGND.n436 VGND.n74 4044.64
R725 VGND.t45 VGND.n74 3942.35
R726 VGND.n444 VGND.n73 3472.59
R727 VGND.n458 VGND.n457 3462.51
R728 VGND.n135 VGND.n134 3164.24
R729 VGND.n137 VGND.n136 3164.24
R730 VGND.n136 VGND.n133 3154.4
R731 VGND.n123 VGND.n122 3108.35
R732 VGND.n126 VGND.n123 3022.83
R733 VGND.n135 VGND.n131 2949.38
R734 VGND.n120 VGND.n76 2758.39
R735 VGND.n444 VGND.n443 2554.5
R736 VGND.n457 VGND.t66 2387.95
R737 VGND.n306 VGND 2380.9
R738 VGND.n145 VGND.n76 2252.33
R739 VGND.n444 VGND.n440 2096.68
R740 VGND.n309 VGND.n308 1953.47
R741 VGND.n459 VGND.n62 1821.62
R742 VGND.n125 VGND.t28 1524.56
R743 VGND.n315 VGND.n77 1397.72
R744 VGND.n305 VGND.t8 1303.08
R745 VGND.n127 VGND.n126 1261.32
R746 VGND.n436 VGND.n435 1170
R747 VGND.n305 VGND.n304 1170
R748 VGND.n451 VGND.n64 1170
R749 VGND.n66 VGND.n63 1170
R750 VGND.n456 VGND.n455 1170
R751 VGND.n443 VGND.n442 1170
R752 VGND.n461 VGND.n460 1170
R753 VGND.n447 VGND.n446 1170
R754 VGND.n379 VGND.n73 1170
R755 VGND.n308 VGND.n307 1170
R756 VGND.n311 VGND.n310 1170
R757 VGND.n143 VGND.n142 1170
R758 VGND.n133 VGND.n132 1170
R759 VGND.n125 VGND.n124 1170
R760 VGND.n483 VGND.n482 1170
R761 VGND.n24 VGND.n2 1170
R762 VGND.n128 VGND.n127 1170
R763 VGND.n489 VGND.n488 1170
R764 VGND.n483 VGND.t34 1134.17
R765 VGND.n309 VGND.n145 1052.01
R766 VGND.t81 VGND.n459 876.702
R767 VGND.n75 VGND.t78 844.357
R768 VGND.n61 VGND.n4 843.24
R769 VGND.t2 VGND.n487 753.322
R770 VGND.n119 VGND.n77 747.253
R771 VGND.t24 VGND.n63 713.466
R772 VGND.t74 VGND.n1 696.106
R773 VGND.n457 VGND.n64 634.212
R774 VGND.t72 VGND.n77 629.832
R775 VGND.n302 VGND.n146 595.942
R776 VGND.n302 VGND.n301 595.942
R777 VGND.n487 VGND.n2 585.742
R778 VGND.n488 VGND.n1 546.058
R779 VGND.t66 VGND.n456 508.485
R780 VGND.n444 VGND.n74 493.118
R781 VGND.n119 VGND.t41 467.337
R782 VGND.t10 VGND.n436 380.034
R783 VGND.n446 VGND.n445 333.548
R784 VGND.n131 VGND.t50 302.156
R785 VGND.n489 VGND.t3 282.339
R786 VGND.n24 VGND.t35 282.339
R787 VGND.n482 VGND.t27 282.339
R788 VGND.n461 VGND.t82 282.339
R789 VGND.n442 VGND.t31 282.339
R790 VGND.n132 VGND.t63 282.339
R791 VGND.n142 VGND.t37 282.339
R792 VGND.n124 VGND.t29 282.339
R793 VGND.n128 VGND.t75 282.339
R794 VGND.n134 VGND.t39 282.339
R795 VGND.n455 VGND.t67 282.339
R796 VGND.n435 VGND.t11 282.339
R797 VGND.n307 VGND.t73 282.339
R798 VGND.n311 VGND.t51 282.339
R799 VGND.n137 VGND.t61 282.339
R800 VGND.n315 VGND.t42 282.339
R801 VGND.n304 VGND.t9 282.339
R802 VGND.n379 VGND.t79 282.339
R803 VGND.n447 VGND.t44 282.339
R804 VGND.n451 VGND.t65 282.339
R805 VGND.n66 VGND.t25 282.339
R806 VGND.t78 VGND.n73 266.457
R807 VGND.n190 VGND.t12 251
R808 VGND.n224 VGND.t17 251
R809 VGND.n281 VGND.t48 251
R810 VGND.t30 VGND.n441 248.936
R811 VGND.n177 VGND.t5 243.028
R812 VGND.n157 VGND.t33 243.028
R813 VGND.n294 VGND.t54 243.028
R814 VGND.n135 VGND.t38 236.923
R815 VGND.n309 VGND.n306 219.505
R816 VGND.n164 VGND.n163 218.506
R817 VGND.n226 VGND.n151 218.506
R818 VGND.n248 VGND.n247 218.506
R819 VGND.n126 VGND.n125 212.281
R820 VGND.n143 VGND.n122 204.773
R821 VGND.n161 VGND.n160 200.201
R822 VGND.n233 VGND.n232 200.201
R823 VGND.n251 VGND.n250 200.201
R824 VGND.n173 VGND.n172 199.739
R825 VGND.n207 VGND.n206 199.739
R826 VGND.n239 VGND.n238 199.739
R827 VGND.n183 VGND.n168 199.53
R828 VGND.n155 VGND.n154 199.53
R829 VGND.n288 VGND.n243 199.53
R830 VGND.n456 VGND.n65 190.542
R831 VGND.n443 VGND.t30 187.446
R832 VGND.n144 VGND.t36 183.096
R833 VGND.n488 VGND.t2 170.459
R834 VGND.n308 VGND.t72 169.868
R835 VGND.t34 VGND.n2 166.094
R836 VGND.n306 VGND.n74 165.339
R837 VGND.n444 VGND.t43 159.488
R838 VGND.n127 VGND.t74 158.115
R839 VGND.n458 VGND.n63 144.5
R840 VGND.t36 VGND.n143 140.434
R841 VGND.n445 VGND.t64 132.02
R842 VGND.t18 VGND.n72 128.904
R843 VGND.n460 VGND.t81 124.144
R844 VGND.n446 VGND.t43 122.326
R845 VGND.t62 VGND.n131 120.314
R846 VGND.n310 VGND.t50 111.326
R847 VGND.n145 VGND.n144 104.849
R848 VGND VGND.t20 102.412
R849 VGND.t64 VGND.n64 101.258
R850 VGND.n484 VGND.n4 100.996
R851 VGND.t4 VGND.n118 94.8614
R852 VGND.t0 VGND.t56 93.0774
R853 VGND.n133 VGND.t62 92.2804
R854 VGND.n168 VGND.t57 74.8666
R855 VGND.n154 VGND.t69 74.8666
R856 VGND.n243 VGND.t77 74.8666
R857 VGND.n136 VGND.t60 55.9751
R858 VGND.n160 VGND.t15 54.2862
R859 VGND.n232 VGND.t16 54.2862
R860 VGND.n250 VGND.t46 54.2862
R861 VGND.n484 VGND.n483 46.6396
R862 VGND VGND.t71 45.7764
R863 VGND.n120 VGND.n3 45.2738
R864 VGND.n460 VGND.n61 40.8576
R865 VGND.n168 VGND.t1 40.0005
R866 VGND.n154 VGND.t40 40.0005
R867 VGND.n243 VGND.t32 40.0005
R868 VGND.n172 VGND.t22 38.5719
R869 VGND.n172 VGND.t70 38.5719
R870 VGND.n206 VGND.t7 38.5719
R871 VGND.n206 VGND.t80 38.5719
R872 VGND.n238 VGND.t53 38.5719
R873 VGND.n238 VGND.t52 38.5719
R874 VGND.n310 VGND.n309 36.639
R875 VGND.n195 VGND.n194 34.6358
R876 VGND.n196 VGND.n195 34.6358
R877 VGND.n185 VGND.n184 34.6358
R878 VGND.n185 VGND.n166 34.6358
R879 VGND.n189 VGND.n166 34.6358
R880 VGND.n178 VGND.n170 34.6358
R881 VGND.n182 VGND.n170 34.6358
R882 VGND.n213 VGND.n212 34.6358
R883 VGND.n214 VGND.n213 34.6358
R884 VGND.n219 VGND.n218 34.6358
R885 VGND.n220 VGND.n219 34.6358
R886 VGND.n220 VGND.n152 34.6358
R887 VGND.n227 VGND.n149 34.6358
R888 VGND.n231 VGND.n149 34.6358
R889 VGND.n293 VGND.n241 34.6358
R890 VGND.n289 VGND.n241 34.6358
R891 VGND.n287 VGND.n244 34.6358
R892 VGND.n283 VGND.n244 34.6358
R893 VGND.n283 VGND.n282 34.6358
R894 VGND.n277 VGND.n276 34.6358
R895 VGND.n276 VGND.n275 34.6358
R896 VGND.n191 VGND.n164 32.7534
R897 VGND.n226 VGND.n225 32.7534
R898 VGND.n280 VGND.n248 32.7534
R899 VGND.n191 VGND.n190 31.2476
R900 VGND.n225 VGND.n224 31.2476
R901 VGND.n281 VGND.n280 31.2476
R902 VGND.n183 VGND.n182 30.8711
R903 VGND.n214 VGND.n155 30.8711
R904 VGND.n289 VGND.n288 30.8711
R905 VGND.n178 VGND.n177 27.4829
R906 VGND.n212 VGND.n157 27.4829
R907 VGND.n294 VGND.n293 27.4829
R908 VGND.t6 VGND.t68 27.1458
R909 VGND.n160 VGND.t49 25.9346
R910 VGND.n232 VGND.t76 25.9346
R911 VGND.n250 VGND.t55 25.9346
R912 VGND.t58 VGND.t0 25.3851
R913 VGND.n163 VGND.t59 24.9236
R914 VGND.n163 VGND.t14 24.9236
R915 VGND.n151 VGND.t23 24.9236
R916 VGND.n151 VGND.t19 24.9236
R917 VGND.n247 VGND.t21 24.9236
R918 VGND.n247 VGND.t47 24.9236
R919 VGND.n201 VGND.n200 23.7181
R920 VGND.n196 VGND.n161 23.7181
R921 VGND.n205 VGND.n159 23.7181
R922 VGND.n233 VGND.n231 23.7181
R923 VGND.n234 VGND.n147 23.7181
R924 VGND.n300 VGND.n299 23.7181
R925 VGND.n275 VGND.n251 23.7181
R926 VGND.n176 VGND.n173 22.9652
R927 VGND.n177 VGND.n176 22.9652
R928 VGND.n208 VGND.n207 22.9652
R929 VGND.n208 VGND.n157 22.9652
R930 VGND.n295 VGND.n239 22.9652
R931 VGND.n295 VGND.n294 22.9652
R932 VGND.n190 VGND.n189 22.2123
R933 VGND.n224 VGND.n152 22.2123
R934 VGND.n282 VGND.n281 22.2123
R935 VGND.n200 VGND.n161 21.4593
R936 VGND.n207 VGND.n205 21.4593
R937 VGND.n234 VGND.n233 21.4593
R938 VGND.n299 VGND.n239 21.4593
R939 VGND.n141 VGND.n130 20.9265
R940 VGND.n131 VGND.n122 20.0607
R941 VGND.t18 VGND.t45 19.8983
R942 VGND.t18 VGND.n302 19.7425
R943 VGND VGND.n272 17.3883
R944 VGND.n463 VGND.n60 17.0502
R945 VGND.n440 VGND.n76 14.7835
R946 VGND.n435 VGND.n434 13.3141
R947 VGND.n307 VGND.n98 13.3141
R948 VGND.n312 VGND.n311 13.3141
R949 VGND.n138 VGND.n137 13.3141
R950 VGND.n316 VGND.n315 13.3141
R951 VGND.n304 VGND.n303 13.3141
R952 VGND.n380 VGND.n379 13.3141
R953 VGND.n448 VGND.n447 13.3141
R954 VGND.n452 VGND.n451 13.3141
R955 VGND.n67 VGND.n66 13.3141
R956 VGND VGND.n24 13.2586
R957 VGND.n482 VGND 13.2586
R958 VGND VGND.n461 13.2586
R959 VGND.n442 VGND 13.2586
R960 VGND.n132 VGND 13.2586
R961 VGND.n142 VGND 13.2586
R962 VGND.n124 VGND 13.2586
R963 VGND VGND.n128 13.2586
R964 VGND.n134 VGND 13.2586
R965 VGND.n455 VGND 13.2586
R966 VGND VGND.n489 13.2586
R967 VGND VGND.n60 10.8878
R968 VGND.n184 VGND.n183 10.5417
R969 VGND.n218 VGND.n155 10.5417
R970 VGND.n288 VGND.n287 10.5417
R971 VGND.n453 VGND.n450 9.52816
R972 VGND VGND.n454 9.46719
R973 VGND.n275 VGND.n274 9.3005
R974 VGND.n276 VGND.n249 9.3005
R975 VGND.n278 VGND.n277 9.3005
R976 VGND.n280 VGND.n279 9.3005
R977 VGND.n281 VGND.n246 9.3005
R978 VGND.n282 VGND.n245 9.3005
R979 VGND.n284 VGND.n283 9.3005
R980 VGND.n285 VGND.n244 9.3005
R981 VGND.n287 VGND.n286 9.3005
R982 VGND.n288 VGND.n242 9.3005
R983 VGND.n290 VGND.n289 9.3005
R984 VGND.n291 VGND.n241 9.3005
R985 VGND.n293 VGND.n292 9.3005
R986 VGND.n294 VGND.n240 9.3005
R987 VGND.n296 VGND.n295 9.3005
R988 VGND.n297 VGND.n239 9.3005
R989 VGND.n299 VGND.n298 9.3005
R990 VGND.n300 VGND.n237 9.3005
R991 VGND.n176 VGND.n175 9.3005
R992 VGND.n177 VGND.n171 9.3005
R993 VGND.n179 VGND.n178 9.3005
R994 VGND.n180 VGND.n170 9.3005
R995 VGND.n182 VGND.n181 9.3005
R996 VGND.n183 VGND.n169 9.3005
R997 VGND.n184 VGND.n167 9.3005
R998 VGND.n186 VGND.n185 9.3005
R999 VGND.n187 VGND.n166 9.3005
R1000 VGND.n189 VGND.n188 9.3005
R1001 VGND.n190 VGND.n165 9.3005
R1002 VGND.n192 VGND.n191 9.3005
R1003 VGND.n194 VGND.n193 9.3005
R1004 VGND.n195 VGND.n162 9.3005
R1005 VGND.n197 VGND.n196 9.3005
R1006 VGND.n198 VGND.n161 9.3005
R1007 VGND.n200 VGND.n199 9.3005
R1008 VGND.n203 VGND.n159 9.3005
R1009 VGND.n205 VGND.n204 9.3005
R1010 VGND.n207 VGND.n158 9.3005
R1011 VGND.n209 VGND.n208 9.3005
R1012 VGND.n210 VGND.n157 9.3005
R1013 VGND.n212 VGND.n211 9.3005
R1014 VGND.n213 VGND.n156 9.3005
R1015 VGND.n215 VGND.n214 9.3005
R1016 VGND.n216 VGND.n155 9.3005
R1017 VGND.n218 VGND.n217 9.3005
R1018 VGND.n219 VGND.n153 9.3005
R1019 VGND.n221 VGND.n220 9.3005
R1020 VGND.n222 VGND.n152 9.3005
R1021 VGND.n224 VGND.n223 9.3005
R1022 VGND.n225 VGND.n150 9.3005
R1023 VGND.n228 VGND.n227 9.3005
R1024 VGND.n229 VGND.n149 9.3005
R1025 VGND.n231 VGND.n230 9.3005
R1026 VGND.n233 VGND.n148 9.3005
R1027 VGND.n235 VGND.n234 9.3005
R1028 VGND.n236 VGND.n147 9.3005
R1029 VGND.n202 VGND.n201 9.3005
R1030 VGND.n139 VGND.n138 9.16992
R1031 VGND VGND.n141 8.69654
R1032 VGND.n313 VGND.n312 8.60727
R1033 VGND.n462 VGND 8.50779
R1034 VGND.n314 VGND.n313 8.47796
R1035 VGND.n68 VGND.n67 7.73586
R1036 VGND.n140 VGND 7.66873
R1037 VGND.t20 VGND.t6 7.40375
R1038 VGND VGND.n481 7.24133
R1039 VGND.n317 VGND.n316 7.18609
R1040 VGND.n174 VGND.n173 7.12576
R1041 VGND.n273 VGND.n251 7.12063
R1042 VGND.n453 VGND.n452 6.8256
R1043 VGND VGND.n117 6.67637
R1044 VGND.n449 VGND.n448 6.61112
R1045 VGND.n336 VGND.n98 6.60276
R1046 VGND.n25 VGND 6.5915
R1047 VGND VGND.n0 6.55995
R1048 VGND.n159 VGND.n146 6.367
R1049 VGND.n301 VGND.n147 6.367
R1050 VGND.n301 VGND.n300 6.367
R1051 VGND.n201 VGND.n146 6.367
R1052 VGND.n130 VGND 6.30778
R1053 VGND.n413 VGND.n380 6.21471
R1054 VGND.n129 VGND 6.20286
R1055 VGND.n303 VGND.n78 6.13644
R1056 VGND.n434 VGND.n433 5.99894
R1057 VGND.n272 VGND.n270 4.82646
R1058 VGND.t56 VGND.t13 4.23127
R1059 VGND.n313 VGND.n117 3.52873
R1060 VGND.n271 VGND 3.40017
R1061 VGND.t71 VGND.t4 3.3096
R1062 VGND.n272 VGND.n271 3.28674
R1063 VGND.n130 VGND.n129 2.92676
R1064 VGND.n454 VGND.n453 2.38171
R1065 VGND.n441 VGND.n65 2.10058
R1066 VGND.n4 VGND.t26 1.91332
R1067 VGND.n194 VGND.n164 1.88285
R1068 VGND.n227 VGND.n226 1.88285
R1069 VGND.n277 VGND.n248 1.88285
R1070 VGND.n141 VGND.n140 1.59945
R1071 VGND.n129 VGND.n0 1.28972
R1072 VGND.t68 VGND.t18 1.23438
R1073 VGND.n271 VGND.n69 1.1273
R1074 VGND.n140 VGND.n139 1.05629
R1075 VGND.n454 VGND.n69 0.953601
R1076 VGND.n139 VGND.n117 0.951859
R1077 VGND.n68 VGND.n60 0.753637
R1078 VGND.n252 uo_out[4] 0.7008
R1079 VGND.n26 VGND.n0 0.663554
R1080 VGND.n359 VGND.n358 0.457033
R1081 VGND.n253 VGND.n252 0.4329
R1082 VGND.n254 VGND.n253 0.4329
R1083 VGND.n255 VGND.n254 0.4329
R1084 VGND.n256 VGND.n255 0.4329
R1085 VGND.n257 VGND.n256 0.4329
R1086 VGND.n258 VGND.n257 0.4329
R1087 VGND.n259 VGND.n258 0.4329
R1088 VGND.n260 VGND.n259 0.4329
R1089 VGND.n261 VGND.n260 0.4329
R1090 VGND.n262 VGND.n261 0.4329
R1091 VGND.n263 VGND.n262 0.4329
R1092 VGND.n264 VGND.n263 0.4329
R1093 VGND.n265 VGND.n264 0.4329
R1094 VGND.n266 VGND.n265 0.4329
R1095 VGND.n267 VGND.n266 0.4329
R1096 VGND.n268 VGND.n267 0.4329
R1097 VGND.n269 VGND.n268 0.4329
R1098 VGND.n270 VGND.n269 0.4329
R1099 VGND.n356 VGND.n78 0.297375
R1100 VGND.n252 uo_out[5] 0.2684
R1101 VGND.n253 uo_out[6] 0.2684
R1102 VGND.n254 uo_out[7] 0.2684
R1103 VGND.n255 uio_out[0] 0.2684
R1104 VGND.n256 uio_out[1] 0.2684
R1105 VGND.n257 uio_out[2] 0.2684
R1106 VGND.n258 uio_out[3] 0.2684
R1107 VGND.n259 uio_out[4] 0.2684
R1108 VGND.n260 uio_out[5] 0.2684
R1109 VGND.n261 uio_out[6] 0.2684
R1110 VGND.n262 uio_out[7] 0.2684
R1111 VGND.n263 uio_oe[0] 0.2684
R1112 VGND.n264 uio_oe[1] 0.2684
R1113 VGND.n265 uio_oe[2] 0.2684
R1114 VGND.n266 uio_oe[3] 0.2684
R1115 VGND.n267 uio_oe[4] 0.2684
R1116 VGND.n268 uio_oe[5] 0.2684
R1117 VGND.n269 uio_oe[6] 0.2684
R1118 VGND.n270 uio_oe[7] 0.2684
R1119 VGND.n356 VGND.n355 0.240747
R1120 VGND.n43 VGND.n7 0.232444
R1121 VGND.n355 VGND.n354 0.201889
R1122 VGND.n354 VGND.n353 0.183192
R1123 VGND.n450 VGND.n70 0.181207
R1124 VGND.n27 VGND.n26 0.177735
R1125 VGND.n317 VGND.n314 0.15732
R1126 VGND.n464 VGND.n463 0.155253
R1127 VGND.n273 VGND 0.152603
R1128 VGND.n44 VGND.n43 0.152388
R1129 VGND.n274 VGND.n273 0.148519
R1130 VGND.n352 VGND.n351 0.145639
R1131 VGND.n413 VGND.n412 0.14536
R1132 VGND.n353 VGND.n352 0.14425
R1133 VGND.n175 VGND.n174 0.143396
R1134 VGND.n355 VGND.n79 0.135917
R1135 VGND.n357 VGND.n356 0.135115
R1136 VGND.n353 VGND.n81 0.134528
R1137 VGND.n354 VGND.n80 0.133742
R1138 VGND.n358 VGND.n78 0.133539
R1139 VGND.n351 VGND.n83 0.133139
R1140 VGND.n352 VGND.n82 0.133139
R1141 VGND.n350 VGND.n84 0.13175
R1142 VGND.n28 VGND.n22 0.131182
R1143 VGND.n347 VGND.n87 0.131118
R1144 VGND.n349 VGND.n85 0.131056
R1145 VGND.n348 VGND.n86 0.130361
R1146 VGND.n343 VGND.n91 0.129761
R1147 VGND.n30 VGND.n20 0.129761
R1148 VGND.n346 VGND.n88 0.129713
R1149 VGND.n27 VGND.n23 0.129713
R1150 VGND.n31 VGND.n19 0.128341
R1151 VGND.n344 VGND.n90 0.128309
R1152 VGND.n29 VGND.n21 0.128309
R1153 VGND.n345 VGND.n89 0.128278
R1154 VGND.n36 VGND.n14 0.12768
R1155 VGND.n34 VGND.n16 0.127655
R1156 VGND.n341 VGND.n93 0.127631
R1157 VGND.n432 VGND.n360 0.127631
R1158 VGND.n32 VGND.n18 0.127631
R1159 VGND.n37 VGND.n13 0.126953
R1160 VGND.n35 VGND.n15 0.126937
R1161 VGND.n340 VGND.n94 0.12692
R1162 VGND.n431 VGND.n361 0.12692
R1163 VGND.n33 VGND.n17 0.12692
R1164 VGND.n342 VGND.n92 0.126904
R1165 VGND.n399 VGND.n394 0.126368
R1166 VGND.n464 VGND.n59 0.126345
R1167 VGND.n466 VGND.n57 0.126333
R1168 VGND.n468 VGND.n55 0.126322
R1169 VGND.n470 VGND.n53 0.126312
R1170 VGND.n42 VGND.n8 0.126244
R1171 VGND.n337 VGND.n97 0.126218
R1172 VGND.n428 VGND.n364 0.126218
R1173 VGND.n339 VGND.n95 0.12621
R1174 VGND.n430 VGND.n362 0.12621
R1175 VGND.n333 VGND.n101 0.1255
R1176 VGND.n334 VGND.n100 0.1255
R1177 VGND.n335 VGND.n99 0.1255
R1178 VGND.n338 VGND.n96 0.1255
R1179 VGND.n429 VGND.n363 0.1255
R1180 VGND.n427 VGND.n365 0.1255
R1181 VGND.n426 VGND.n366 0.1255
R1182 VGND.n425 VGND.n367 0.1255
R1183 VGND.n38 VGND.n12 0.1255
R1184 VGND.n39 VGND.n11 0.1255
R1185 VGND.n40 VGND.n10 0.1255
R1186 VGND.n475 VGND.n48 0.1255
R1187 VGND.n473 VGND.n50 0.1255
R1188 VGND.n465 VGND.n58 0.1255
R1189 VGND.n330 VGND.n104 0.124765
R1190 VGND.n422 VGND.n370 0.124765
R1191 VGND.n41 VGND.n9 0.124765
R1192 VGND.n481 VGND.n480 0.124747
R1193 VGND.n478 VGND.n45 0.124738
R1194 VGND.n476 VGND.n47 0.124728
R1195 VGND.n472 VGND.n51 0.124709
R1196 VGND.n407 VGND.n386 0.124688
R1197 VGND.n405 VGND.n388 0.124678
R1198 VGND.n403 VGND.n390 0.124667
R1199 VGND.n401 VGND.n392 0.124655
R1200 VGND.n400 VGND.n393 0.124655
R1201 VGND.n398 VGND.n395 0.124644
R1202 VGND.n332 VGND.n102 0.124047
R1203 VGND.n424 VGND.n368 0.124047
R1204 VGND.n328 VGND.n106 0.124012
R1205 VGND.n420 VGND.n372 0.124012
R1206 VGND.n326 VGND.n108 0.123994
R1207 VGND.n418 VGND.n374 0.123994
R1208 VGND.n479 VGND.n6 0.123994
R1209 VGND.n477 VGND.n46 0.123976
R1210 VGND.n320 VGND.n114 0.123938
R1211 VGND.n318 VGND.n116 0.123918
R1212 VGND.n410 VGND.n383 0.123918
R1213 VGND.n471 VGND.n52 0.123918
R1214 VGND.n469 VGND.n54 0.123897
R1215 VGND.n467 VGND.n56 0.123877
R1216 VGND.n402 VGND.n391 0.123833
R1217 VGND.n412 VGND.n411 0.123779
R1218 VGND.n331 VGND.n103 0.12332
R1219 VGND.n423 VGND.n369 0.12332
R1220 VGND.n329 VGND.n105 0.123294
R1221 VGND.n421 VGND.n371 0.123294
R1222 VGND.n327 VGND.n107 0.123268
R1223 VGND.n419 VGND.n373 0.123268
R1224 VGND.n325 VGND.n109 0.123241
R1225 VGND.n417 VGND.n375 0.123241
R1226 VGND.n323 VGND.n111 0.123213
R1227 VGND.n321 VGND.n113 0.123185
R1228 VGND.n474 VGND.n49 0.123185
R1229 VGND.n409 VGND.n384 0.123127
R1230 VGND.n324 VGND.n110 0.122488
R1231 VGND.n416 VGND.n376 0.122488
R1232 VGND.n322 VGND.n112 0.122451
R1233 VGND.n408 VGND.n385 0.122335
R1234 VGND.n406 VGND.n387 0.122295
R1235 VGND.n404 VGND.n389 0.122253
R1236 VGND.n319 VGND.n115 0.121642
R1237 VGND.n411 VGND.n382 0.121642
R1238 VGND.n351 VGND.n350 0.120386
R1239 VGND.n175 VGND.n171 0.120292
R1240 VGND.n179 VGND.n171 0.120292
R1241 VGND.n180 VGND.n179 0.120292
R1242 VGND.n181 VGND.n180 0.120292
R1243 VGND.n181 VGND.n169 0.120292
R1244 VGND.n169 VGND.n167 0.120292
R1245 VGND.n186 VGND.n167 0.120292
R1246 VGND.n187 VGND.n186 0.120292
R1247 VGND.n188 VGND.n187 0.120292
R1248 VGND.n188 VGND.n165 0.120292
R1249 VGND.n192 VGND.n165 0.120292
R1250 VGND.n193 VGND.n192 0.120292
R1251 VGND.n193 VGND.n162 0.120292
R1252 VGND.n197 VGND.n162 0.120292
R1253 VGND.n198 VGND.n197 0.120292
R1254 VGND.n199 VGND.n198 0.120292
R1255 VGND.n209 VGND.n158 0.120292
R1256 VGND.n210 VGND.n209 0.120292
R1257 VGND.n211 VGND.n210 0.120292
R1258 VGND.n211 VGND.n156 0.120292
R1259 VGND.n215 VGND.n156 0.120292
R1260 VGND.n216 VGND.n215 0.120292
R1261 VGND.n217 VGND.n216 0.120292
R1262 VGND.n217 VGND.n153 0.120292
R1263 VGND.n221 VGND.n153 0.120292
R1264 VGND.n222 VGND.n221 0.120292
R1265 VGND.n223 VGND.n222 0.120292
R1266 VGND.n223 VGND.n150 0.120292
R1267 VGND.n228 VGND.n150 0.120292
R1268 VGND.n229 VGND.n228 0.120292
R1269 VGND.n230 VGND.n229 0.120292
R1270 VGND.n230 VGND.n148 0.120292
R1271 VGND.n235 VGND.n148 0.120292
R1272 VGND.n297 VGND.n296 0.120292
R1273 VGND.n296 VGND.n240 0.120292
R1274 VGND.n292 VGND.n240 0.120292
R1275 VGND.n292 VGND.n291 0.120292
R1276 VGND.n291 VGND.n290 0.120292
R1277 VGND.n290 VGND.n242 0.120292
R1278 VGND.n286 VGND.n242 0.120292
R1279 VGND.n286 VGND.n285 0.120292
R1280 VGND.n285 VGND.n284 0.120292
R1281 VGND.n284 VGND.n245 0.120292
R1282 VGND.n246 VGND.n245 0.120292
R1283 VGND.n279 VGND.n246 0.120292
R1284 VGND.n279 VGND.n278 0.120292
R1285 VGND.n278 VGND.n249 0.120292
R1286 VGND.n274 VGND.n249 0.120292
R1287 VGND.n397 VGND.n71 0.115369
R1288 VGND.n350 VGND.n349 0.112306
R1289 VGND.n399 VGND.n398 0.111879
R1290 VGND.n398 VGND.n397 0.111186
R1291 VGND.n349 VGND.n348 0.109795
R1292 VGND.n401 VGND.n400 0.108943
R1293 VGND.n43 VGND.n42 0.108833
R1294 VGND.n400 VGND.n399 0.107764
R1295 VGND.n348 VGND.n347 0.107742
R1296 VGND.n402 VGND.n401 0.107535
R1297 VGND.n314 VGND.n116 0.107341
R1298 VGND.n403 VGND.n402 0.106725
R1299 VGND.n465 VGND.n464 0.106074
R1300 VGND.n466 VGND.n465 0.105969
R1301 VGND.n405 VGND.n404 0.1059
R1302 VGND.n467 VGND.n466 0.105163
R1303 VGND.n404 VGND.n403 0.104834
R1304 VGND.n406 VGND.n405 0.104121
R1305 VGND.n407 VGND.n406 0.103867
R1306 VGND.n468 VGND.n467 0.10332
R1307 VGND.n469 VGND.n468 0.10304
R1308 VGND.n29 VGND.n28 0.102984
R1309 VGND.n471 VGND.n470 0.102502
R1310 VGND.n410 VGND.n409 0.102274
R1311 VGND.n408 VGND.n407 0.10217
R1312 VGND.n409 VGND.n408 0.101442
R1313 VGND.n470 VGND.n469 0.101279
R1314 VGND.n320 VGND.n319 0.1005
R1315 VGND.n473 VGND.n472 0.100144
R1316 VGND.n321 VGND.n320 0.0994435
R1317 VGND.n474 VGND.n473 0.099433
R1318 VGND.n472 VGND.n471 0.0992982
R1319 VGND.n319 VGND.n318 0.0991552
R1320 VGND.n411 VGND.n410 0.0991552
R1321 VGND VGND.n158 0.0981562
R1322 VGND VGND.n297 0.0981562
R1323 VGND.n381 VGND.n378 0.0981562
R1324 VGND.n323 VGND.n322 0.0977932
R1325 VGND.n415 VGND.n414 0.0977932
R1326 VGND.n476 VGND.n475 0.0976284
R1327 VGND.n324 VGND.n323 0.0968228
R1328 VGND.n416 VGND.n415 0.0968228
R1329 VGND.n322 VGND.n321 0.0966929
R1330 VGND.n477 VGND.n476 0.0965648
R1331 VGND.n475 VGND.n474 0.0962384
R1332 VGND.n325 VGND.n324 0.0962186
R1333 VGND.n417 VGND.n416 0.0962186
R1334 VGND.n394 VGND.n393 0.0959861
R1335 VGND.n326 VGND.n325 0.0956231
R1336 VGND.n418 VGND.n417 0.0956231
R1337 VGND.n478 VGND.n477 0.0955348
R1338 VGND.n479 VGND.n478 0.0948777
R1339 VGND.n395 VGND.n394 0.0946781
R1340 VGND.n31 VGND.n30 0.0945657
R1341 VGND.n28 VGND.n27 0.0938949
R1342 VGND.n346 VGND.n345 0.0937672
R1343 VGND.n30 VGND.n29 0.0931452
R1344 VGND.n344 VGND.n343 0.0930016
R1345 VGND.n415 VGND.n377 0.0927256
R1346 VGND.n327 VGND.n326 0.0927181
R1347 VGND.n419 VGND.n418 0.0927181
R1348 VGND.n347 VGND.n346 0.0923627
R1349 VGND.n7 VGND.n5 0.0921667
R1350 VGND.n328 VGND.n327 0.0920855
R1351 VGND.n420 VGND.n419 0.0920855
R1352 VGND.n480 VGND.n479 0.0919467
R1353 VGND.n345 VGND.n344 0.0914722
R1354 VGND.n480 VGND.n44 0.0912494
R1355 VGND.n329 VGND.n328 0.091171
R1356 VGND.n421 VGND.n420 0.091171
R1357 VGND.n32 VGND.n31 0.0904148
R1358 VGND.n392 VGND.n391 0.090027
R1359 VGND.n393 VGND.n392 0.090027
R1360 VGND.n330 VGND.n329 0.0898264
R1361 VGND.n422 VGND.n421 0.0898264
R1362 VGND.n332 VGND.n331 0.0891127
R1363 VGND.n424 VGND.n423 0.0891127
R1364 VGND.n38 VGND.n37 0.0881565
R1365 VGND.n42 VGND.n41 0.0881488
R1366 VGND.n41 VGND.n40 0.0879493
R1367 VGND.n333 VGND.n332 0.0878131
R1368 VGND.n425 VGND.n424 0.0878131
R1369 VGND.n331 VGND.n330 0.0876124
R1370 VGND.n423 VGND.n422 0.0876124
R1371 VGND.n33 VGND.n32 0.0875536
R1372 VGND.n391 VGND.n390 0.0871667
R1373 VGND.n37 VGND.n36 0.0868953
R1374 VGND.n462 VGND.n59 0.0866486
R1375 VGND.n36 VGND.n35 0.0863769
R1376 VGND.n342 VGND.n341 0.0859735
R1377 VGND.n35 VGND.n34 0.0856762
R1378 VGND.n44 VGND.n5 0.085541
R1379 VGND.n390 VGND.n389 0.0855
R1380 VGND.n34 VGND.n33 0.0852048
R1381 VGND.n343 VGND.n342 0.0851591
R1382 VGND.n40 VGND.n39 0.0850588
R1383 VGND.n59 VGND.n58 0.0838333
R1384 VGND.n341 VGND.n340 0.0835966
R1385 VGND.n432 VGND.n431 0.0835966
R1386 VGND.n428 VGND.n427 0.0833636
R1387 VGND.n334 VGND.n333 0.0833488
R1388 VGND.n426 VGND.n425 0.0833488
R1389 VGND.n39 VGND.n38 0.0833488
R1390 VGND.n429 VGND.n428 0.0825455
R1391 VGND.n58 VGND.n57 0.0821667
R1392 VGND.n336 VGND.n335 0.081981
R1393 VGND.n339 VGND.n338 0.0819394
R1394 VGND.n430 VGND.n429 0.0819394
R1395 VGND.n335 VGND.n334 0.0816782
R1396 VGND.n427 VGND.n426 0.0816782
R1397 VGND.n389 VGND.n388 0.0816688
R1398 VGND.n340 VGND.n339 0.0813424
R1399 VGND.n431 VGND.n430 0.0813424
R1400 VGND.n388 VGND.n387 0.0810921
R1401 VGND.n412 VGND.n381 0.0797137
R1402 VGND.n449 VGND.n71 0.0796453
R1403 VGND.n396 VGND.n395 0.0796157
R1404 VGND.n57 VGND.n56 0.0784221
R1405 VGND.n56 VGND.n55 0.0778026
R1406 VGND.n387 VGND.n386 0.0774231
R1407 VGND.n386 VGND.n385 0.0767987
R1408 VGND.n397 VGND.n396 0.0762042
R1409 VGND.n174 VGND 0.0758148
R1410 VGND.n55 VGND.n54 0.074218
R1411 VGND.n54 VGND.n53 0.073552
R1412 VGND.n385 VGND.n384 0.0732848
R1413 VGND.n433 VGND.n359 0.0732142
R1414 VGND.n433 VGND.n432 0.0719286
R1415 VGND.n384 VGND.n383 0.0717025
R1416 VGND.n116 VGND.n115 0.0701203
R1417 VGND.n383 VGND.n382 0.0701203
R1418 VGND.n53 VGND.n52 0.0701203
R1419 VGND.n52 VGND.n51 0.068538
R1420 VGND.n51 VGND.n50 0.0669557
R1421 VGND.n115 VGND.n114 0.066858
R1422 VGND.n382 VGND.n381 0.066858
R1423 VGND.n377 VGND.n376 0.0667809
R1424 VGND.n114 VGND.n113 0.066125
R1425 VGND.n113 VGND.n112 0.0637716
R1426 VGND.n50 VGND.n49 0.0637716
R1427 VGND.n49 VGND.n48 0.063
R1428 VGND.n112 VGND.n111 0.0614756
R1429 VGND.n338 VGND.n337 0.0609482
R1430 VGND.n48 VGND.n47 0.0606852
R1431 VGND.n199 VGND 0.0603958
R1432 VGND.n202 VGND 0.0603958
R1433 VGND.n203 VGND 0.0603958
R1434 VGND.n204 VGND 0.0603958
R1435 VGND VGND.n235 0.0603958
R1436 VGND.n236 VGND 0.0603958
R1437 VGND.n237 VGND 0.0603958
R1438 VGND.n298 VGND 0.0603958
R1439 VGND.n111 VGND.n110 0.0599512
R1440 VGND.n47 VGND.n46 0.0584268
R1441 VGND.n110 VGND.n109 0.0577289
R1442 VGND.n376 VGND.n375 0.0577289
R1443 VGND.n46 VGND.n45 0.0569024
R1444 VGND.n109 VGND.n108 0.0562229
R1445 VGND.n375 VGND.n374 0.0562229
R1446 VGND.n434 VGND 0.0560556
R1447 VGND.n98 VGND 0.0560556
R1448 VGND.n312 VGND 0.0560556
R1449 VGND.n138 VGND 0.0560556
R1450 VGND.n316 VGND 0.0560556
R1451 VGND.n303 VGND 0.0560556
R1452 VGND.n380 VGND 0.0560556
R1453 VGND.n448 VGND 0.0560556
R1454 VGND.n452 VGND 0.0560556
R1455 VGND.n67 VGND 0.0560556
R1456 VGND.n450 VGND.n449 0.0554302
R1457 VGND.n108 VGND.n107 0.0547169
R1458 VGND.n374 VGND.n373 0.0547169
R1459 VGND.n45 VGND.n6 0.0547169
R1460 VGND.n481 VGND.n6 0.0532108
R1461 VGND.n107 VGND.n106 0.0525833
R1462 VGND.n373 VGND.n372 0.0525833
R1463 VGND.n396 VGND.n70 0.0514752
R1464 VGND.n106 VGND.n105 0.0510952
R1465 VGND.n372 VGND.n371 0.0510952
R1466 VGND.n105 VGND.n104 0.0490294
R1467 VGND.n371 VGND.n370 0.0490294
R1468 VGND.n360 VGND.n359 0.0488306
R1469 VGND.n8 VGND.n7 0.046631
R1470 VGND.n414 VGND.n378 0.0461288
R1471 VGND.n104 VGND.n103 0.0460882
R1472 VGND.n370 VGND.n369 0.0460882
R1473 VGND.n9 VGND.n8 0.0460882
R1474 VGND.n103 VGND.n102 0.0455581
R1475 VGND.n369 VGND.n368 0.0455581
R1476 VGND.n10 VGND.n9 0.0446176
R1477 VGND.n102 VGND.n101 0.0441047
R1478 VGND.n368 VGND.n367 0.0441047
R1479 VGND.n101 VGND.n100 0.0411977
R1480 VGND.n100 VGND.n99 0.0411977
R1481 VGND.n366 VGND.n365 0.0411977
R1482 VGND.n367 VGND.n366 0.0411977
R1483 VGND.n12 VGND.n11 0.0411977
R1484 VGND.n11 VGND.n10 0.0411977
R1485 VGND.n463 VGND.n462 0.0401474
R1486 VGND.n13 VGND.n12 0.0382907
R1487 VGND.n71 VGND.n70 0.0381773
R1488 VGND.n99 VGND.n97 0.0378563
R1489 VGND.n365 VGND.n364 0.0378563
R1490 VGND.n14 VGND.n13 0.0368372
R1491 VGND.n97 VGND.n96 0.0364195
R1492 VGND.n364 VGND.n363 0.0364195
R1493 VGND.n481 VGND.n5 0.0353361
R1494 VGND.n318 VGND.n317 0.0353101
R1495 VGND.n15 VGND.n14 0.0349828
R1496 VGND.n96 VGND.n95 0.0345909
R1497 VGND.n363 VGND.n362 0.0345909
R1498 VGND VGND.n202 0.0343542
R1499 VGND VGND.n203 0.0343542
R1500 VGND VGND.n236 0.0343542
R1501 VGND VGND.n237 0.0343542
R1502 VGND.n16 VGND.n15 0.033546
R1503 VGND.n95 VGND.n94 0.0331705
R1504 VGND.n362 VGND.n361 0.0331705
R1505 VGND.n94 VGND.n93 0.03175
R1506 VGND.n361 VGND.n360 0.03175
R1507 VGND.n17 VGND.n16 0.03175
R1508 VGND.n378 VGND.n377 0.0315583
R1509 VGND.n93 VGND.n92 0.0303295
R1510 VGND.n18 VGND.n17 0.0303295
R1511 VGND.n19 VGND.n18 0.0289091
R1512 VGND.n92 VGND.n91 0.0285899
R1513 VGND.n91 VGND.n90 0.0260682
R1514 VGND.n20 VGND.n19 0.0260682
R1515 VGND.n90 VGND.n89 0.0257809
R1516 VGND.n21 VGND.n20 0.0257809
R1517 VGND.n22 VGND.n21 0.0232273
R1518 VGND.n88 VGND.n87 0.0229719
R1519 VGND.n23 VGND.n22 0.0229719
R1520 VGND.n89 VGND.n88 0.0227222
R1521 VGND.n204 VGND 0.0226354
R1522 VGND.n298 VGND 0.0226354
R1523 VGND.n87 VGND.n86 0.0201629
R1524 VGND.n25 VGND.n23 0.0199444
R1525 VGND.n86 VGND.n85 0.0185556
R1526 VGND.n85 VGND.n84 0.0171667
R1527 VGND.n69 VGND.n68 0.0169225
R1528 VGND.n414 VGND.n413 0.0158374
R1529 VGND.n84 VGND.n83 0.0157778
R1530 VGND.n83 VGND.n82 0.013
R1531 VGND.n82 VGND.n81 0.013
R1532 VGND.n81 VGND.n80 0.0102222
R1533 VGND.n26 VGND.n25 0.00911038
R1534 VGND.n80 VGND.n79 0.00874176
R1535 VGND.n358 VGND.n357 0.00816087
R1536 VGND.n357 VGND.n79 0.00744444
R1537 VGND.n337 VGND.n336 0.00285443
R1538 uo_out[0] uo_out[0].t0 984.356
R1539 uo_out[0].n0 uo_out[0].t2 582.378
R1540 uo_out[0].n1 uo_out[0].t3 566.953
R1541 uo_out[0].n8 uo_out[0].t1 478.87
R1542 uo_out[0].n1 uo_out[0].n0 424.161
R1543 uo_out[0].n3 uo_out[0].t4 294.557
R1544 uo_out[0].n3 uo_out[0].t5 211.01
R1545 uo_out[0].n2 uo_out[0].n0 204.481
R1546 uo_out[0] uo_out[0].n1 201.921
R1547 uo_out[0].n4 uo_out[0].n3 152
R1548 uo_out[0].n7 uo_out[0].n6 18.3079
R1549 uo_out[0].n5 uo_out[0].n4 17.6405
R1550 uo_out[0].n2 uo_out[0] 10.2405
R1551 uo_out[0] uo_out[0].n8 10.2405
R1552 uo_out[0].n8 uo_out[0].n7 7.5409
R1553 uo_out[0].n6 uo_out[0].n5 6.83545
R1554 uo_out[0].n7 uo_out[0].n2 5.01603
R1555 uo_out[0].n4 uo_out[0] 2.01193
R1556 uo_out[0].n6 uo_out[0] 1.31337
R1557 uo_out[0].n5 uo_out[0] 0.0793043
R1558 uo_out[1].n2 uo_out[1].t0 313.104
R1559 uo_out[1].n0 uo_out[1].t2 294.557
R1560 uo_out[1].t1 uo_out[1].n2 265.769
R1561 uo_out[1] uo_out[1].t1 262.318
R1562 uo_out[1].n0 uo_out[1].t3 211.01
R1563 uo_out[1].n1 uo_out[1].n0 152
R1564 uo_out[1].n5 uo_out[1] 12.6752
R1565 uo_out[1].n4 uo_out[1].n1 11.6411
R1566 uo_out[1].n4 uo_out[1].n3 9.3005
R1567 uo_out[1].n3 uo_out[1] 7.17626
R1568 uo_out[1].n3 uo_out[1].n2 4.84898
R1569 uo_out[1].n5 uo_out[1].n4 4.5029
R1570 uo_out[1].n1 uo_out[1] 1.37896
R1571 uo_out[1] uo_out[1].n5 0.0730806
R1572 uo_out[3].n0 uo_out[3].t0 313.104
R1573 uo_out[3].t1 uo_out[3].n0 265.769
R1574 uo_out[3] uo_out[3].t1 262.318
R1575 uo_out[3].n2 uo_out[3] 19.5328
R1576 uo_out[3].n2 uo_out[3].n1 13.8005
R1577 uo_out[3].n1 uo_out[3].n0 7.17626
R1578 uo_out[3].n1 uo_out[3] 4.84898
R1579 uo_out[3] uo_out[3].n2 0.0529194
C0 m3_10514_15880# m4_10514_15880# 65.3249f
C1 m2_12074_25760# m3_12074_25760# 98.466896f
C2 m1_10514_15880# m2_10514_15880# 0.104063p
C3 m2_12074_25760# m1_12074_25760# 0.152927p
C4 m3_10514_15880# m2_10514_15880# 67.004105f
C5 m4_12074_25760# m3_12074_25760# 95.99921f
C6 uo_out[0] VGND 9.161079f
C7 uo_out[3] VGND 1.95825f
C8 VPWR VGND 0.161567p
C9 m4_10514_15880# VGND 11.0708f $ **FLOATING
C10 m4_12074_25760# VGND 8.74739f $ **FLOATING
C11 m3_10514_15880# VGND 12.571401f $ **FLOATING
C12 m3_12074_25760# VGND 10.2012f $ **FLOATING
C13 m2_10514_15880# VGND 11.5358f $ **FLOATING
C14 m2_12074_25760# VGND 9.56448f $ **FLOATING
C15 m1_10514_15880# VGND 32.9027f $ **FLOATING
C16 m1_12074_25760# VGND 40.2807f $ **FLOATING
C17 ring_0/skullfet_inverter_16.A VGND 4.53396f
C18 ring_0/skullfet_inverter_17.A VGND 4.70918f
C19 ring_0/skullfet_inverter_15.A VGND 4.82841f
C20 ring_0/skullfet_inverter_18.A VGND 4.90629f
C21 ring_0/skullfet_inverter_14.A VGND 4.98419f
C22 ring_0/skullfet_inverter_19.A VGND 4.923029f
C23 ring_0/skullfet_inverter_13.A VGND 4.78946f
C24 ring_0/skullfet_inverter_20.A VGND 4.72064f
C25 ring_0/skullfet_inverter_12.A VGND 5.60339f
C26 ring_0/skullfet_inverter_20.Y VGND 5.35745f
C27 ring_0/skullfet_inverter_11.A VGND 4.97718f
C28 ring_0/skullfet_inverter_1.A VGND 5.16765f
C29 ring_0/skullfet_inverter_10.A VGND 5.58737f
C30 ring_0/skullfet_inverter_2.A VGND 5.65285f
C31 ring_0/skullfet_inverter_9.A VGND 4.78733f
C32 ring_0/skullfet_inverter_3.A VGND 4.92041f
C33 ring_0/skullfet_inverter_4.A VGND 4.93544f
C34 ring_0/skullfet_inverter_8.A VGND 4.94116f
C35 ring_0/skullfet_inverter_7.A VGND 4.81796f
C36 ring_0/skullfet_inverter_6.A VGND 4.53217f
.ends

