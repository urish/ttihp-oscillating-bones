* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] VAPWR
+ VDPWR VGND
X0 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VAPWR.t27 VAPWR.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X1 VGND.t66 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_5.A VGND.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X2 VDPWR.t63 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_10715_43723# VDPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X3 a_10544_44089# a_10297_43723# VDPWR.t57 VDPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X4 a_10297_43723# a_10168_43997# a_9876_43697# VGND.t36 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5 a_10368_43697# a_10161_43697# a_10544_44089# VDPWR.t61 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X6 VGND.t83 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X7 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VAPWR.t31 VAPWR.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X8 VGND.t62 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X9 a_13468_43697# a_13740_43697# VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VDPWR.t17 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12647_43723# VDPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X11 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VAPWR.t33 VAPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X12 VGND.t55 a_11441_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t54 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VAPWR.t23 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VAPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X14 a_12093_43697# uo_out[1].t2 VDPWR.t13 VDPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_12051_44089# a_11536_43697# VDPWR.t37 VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X16 VAPWR.t21 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VAPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X17 a_14232_43697# a_14032_43997# a_14381_43723# VGND.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X18 VGND.t3 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X19 VGND.t69 a_13468_43697# uo_out[1].t0 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 VDPWR.t65 a_9509_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VDPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X21 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VGND.t51 VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X22 ring_0/skullfet_inverter_9.A skullfet_level_shifter.A VAPWR.t7 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X23 a_13960_43723# a_13468_43697# VGND.t68 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t87 VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X25 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t89 VGND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X26 VGND.t95 a_9604_43697# uo_out[3].t0 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t24 VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X28 VAPWR.t41 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VAPWR.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X29 VGND.t5 a_14232_43697# a_14161_43723# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X30 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VAPWR.t35 VAPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X31 VGND.t16 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X32 VGND.t81 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X33 a_12647_43723# a_12100_43997# a_12300_43697# VDPWR.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X34 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t49 VGND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X35 a_13468_43697# a_13740_43697# VDPWR.t45 VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X36 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VAPWR.t11 VAPWR.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X37 a_11441_43697# a_11536_43697# VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X38 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t60 VGND.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X39 VDPWR.t60 a_10161_43697# a_10168_43997# VDPWR.t59 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X40 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_5.A VAPWR.t17 VAPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X41 uo_out[0].t0 skullfet_level_shifter.A VGND.t14 VGND.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X42 a_14025_43697# uo_out[0].t2 VGND.t31 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 a_14232_43697# a_14025_43697# a_14408_44089# VDPWR.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X44 a_14161_43723# a_14025_43697# a_13740_43697# VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 VDPWR.t55 a_13468_43697# uo_out[1].t1 VDPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X46 VDPWR.t41 a_12093_43697# a_12100_43997# VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X47 VDPWR.t71 a_9604_43697# uo_out[3].t1 VDPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X48 VGND.t30 a_14025_43697# a_14032_43997# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X49 a_9509_43697# a_9604_43697# VDPWR.t69 VDPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X50 VGND.t1 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X51 a_10119_44089# a_9604_43697# VDPWR.t67 VDPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X52 a_10161_43697# uo_out[2].t2 VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X53 a_13740_43697# a_14032_43997# a_13983_44089# VDPWR.t3 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X54 VAPWR.t19 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VAPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X55 VGND.t21 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X56 a_12028_43723# a_11536_43697# VGND.t45 VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X57 skullfet_level_shifter.A ring_0/skullfet_inverter_7.A VAPWR.t15 VAPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X58 a_10517_43723# a_10297_43723# VGND.t71 VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X59 VAPWR.t13 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VAPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X60 VGND.t33 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_6.A VGND.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X61 a_9604_43697# a_9876_43697# VGND.t64 VGND.t63 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X62 VGND.t58 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_14579_43723# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X63 a_12093_43697# uo_out[1].t3 VGND.t22 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X64 VAPWR.t25 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VAPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X65 a_12449_43723# a_12229_43723# VGND.t17 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X66 VGND.t43 a_11536_43697# uo_out[2].t0 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X67 VGND.t85 a_9509_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VGND.t77 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X69 VGND.t37 a_12300_43697# a_12229_43723# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X70 a_10715_43723# a_10168_43997# a_10368_43697# VDPWR.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X71 a_9604_43697# a_9876_43697# VDPWR.t49 VDPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X72 a_11536_43697# a_11808_43697# VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X73 a_13373_43697# a_13468_43697# VGND.t67 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X74 a_14408_44089# a_14161_43723# VDPWR.t5 VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X75 VGND.t27 ring_0/skullfet_inverter_7.A skullfet_level_shifter.A VGND.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X76 VGND.t75 a_10161_43697# a_10168_43997# VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X77 a_10096_43723# a_9604_43697# VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X78 VDPWR.t33 a_11536_43697# uo_out[2].t1 VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X79 VDPWR.t73 a_13373_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X80 VDPWR.t47 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_14579_43723# VDPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X81 VGND.t47 a_12093_43697# a_12100_43997# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X82 a_14579_43723# a_14025_43697# a_14232_43697# VGND.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X83 a_14161_43723# a_14032_43997# a_13740_43697# VGND.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X84 a_11808_43697# a_12100_43997# a_12051_44089# VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X85 VAPWR.t39 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VAPWR.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X86 a_10161_43697# uo_out[2].t3 VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X87 VAPWR.t37 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VAPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X88 a_10368_43697# a_10168_43997# a_10517_43723# VGND.t35 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X89 a_11536_43697# a_11808_43697# VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X90 VGND.t39 a_10368_43697# a_10297_43723# VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X91 a_12300_43697# a_12100_43997# a_12449_43723# VGND.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X92 a_11808_43697# a_12093_43697# a_12028_43723# VGND.t46 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X93 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VAPWR.t5 VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X94 VDPWR.t7 skullfet_level_shifter.A uo_out[0].t1 VDPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X95 a_13373_43697# a_13468_43697# VDPWR.t53 VDPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X96 VDPWR.t1 a_14232_43697# a_14161_43723# VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X97 a_13740_43697# a_14025_43697# a_13960_43723# VGND.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X98 a_10297_43723# a_10161_43697# a_9876_43697# VDPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 a_11441_43697# a_11536_43697# VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X100 a_12476_44089# a_12229_43723# VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X101 a_12229_43723# a_12100_43997# a_11808_43697# VGND.t34 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X102 a_12229_43723# a_12093_43697# a_11808_43697# VDPWR.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X103 a_12300_43697# a_12093_43697# a_12476_44089# VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X104 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VAPWR.t9 VAPWR.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X105 a_10715_43723# a_10161_43697# a_10368_43697# VGND.t73 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X106 VDPWR.t43 a_11441_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X107 VGND.t8 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X108 VGND.t12 skullfet_level_shifter.A ring_0/skullfet_inverter_9.A VGND.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X109 VGND.t98 a_13373_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X110 a_9509_43697# a_9604_43697# VGND.t91 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X111 VGND.t79 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_10715_43723# VGND.t78 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X112 a_12647_43723# a_12093_43697# a_12300_43697# VGND.t6 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X113 a_9876_43697# a_10168_43997# a_10119_44089# VDPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X114 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_4.A VAPWR.t29 VAPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X115 a_14381_43723# a_14161_43723# VGND.t10 VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X116 VGND.t25 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12647_43723# VGND.t9 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X117 a_14579_43723# a_14032_43997# a_14232_43697# VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X118 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VGND.t53 VGND.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X119 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X120 VDPWR.t31 a_10368_43697# a_10297_43723# VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X121 a_9876_43697# a_10161_43697# a_10096_43723# VGND.t72 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X122 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VAPWR.t3 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X123 a_14025_43697# uo_out[0].t3 VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X124 a_13983_44089# a_13468_43697# VDPWR.t51 VDPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X125 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t97 VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X126 VDPWR.t29 a_12300_43697# a_12229_43723# VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X127 VDPWR.t21 a_14025_43697# a_14032_43997# VDPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
R0 VAPWR.n52 VAPWR.t19 738.799
R1 VAPWR.n54 VAPWR.t35 738.799
R2 VAPWR.n38 VAPWR.t23 738.799
R3 VAPWR.n34 VAPWR.t21 738.799
R4 VAPWR.n6 VAPWR.t11 738.799
R5 VAPWR.n41 VAPWR.t13 738.799
R6 VAPWR.n44 VAPWR.t39 738.799
R7 VAPWR.n47 VAPWR.t37 738.799
R8 VAPWR.n4 VAPWR.t25 738.799
R9 VAPWR.n2 VAPWR.t41 738.799
R10 VAPWR.n60 VAPWR.t1 738.799
R11 VAPWR.n57 VAPWR.t9 738.799
R12 VAPWR.n32 VAPWR.t5 738.799
R13 VAPWR.n7 VAPWR.t33 738.799
R14 VAPWR.n11 VAPWR.t17 738.799
R15 VAPWR.n22 VAPWR.t27 738.799
R16 VAPWR.n19 VAPWR.t15 738.799
R17 VAPWR.n16 VAPWR.t7 738.799
R18 VAPWR.n13 VAPWR.t3 738.799
R19 VAPWR.n9 VAPWR.t29 738.799
R20 VAPWR.n27 VAPWR.t31 738.799
R21 VAPWR.n60 VAPWR.t0 707.519
R22 VAPWR.n57 VAPWR.t8 707.519
R23 VAPWR.n52 VAPWR.t18 707.519
R24 VAPWR.n54 VAPWR.t34 707.519
R25 VAPWR.n38 VAPWR.t22 707.519
R26 VAPWR.n34 VAPWR.t20 707.519
R27 VAPWR.n32 VAPWR.t4 707.519
R28 VAPWR.n6 VAPWR.t10 707.519
R29 VAPWR.n7 VAPWR.t32 707.519
R30 VAPWR.n11 VAPWR.t16 707.519
R31 VAPWR.n22 VAPWR.t26 707.519
R32 VAPWR.n19 VAPWR.t14 707.519
R33 VAPWR.n16 VAPWR.t6 707.519
R34 VAPWR.n13 VAPWR.t2 707.519
R35 VAPWR.n9 VAPWR.t28 707.519
R36 VAPWR.n27 VAPWR.t30 707.519
R37 VAPWR.n41 VAPWR.t12 707.519
R38 VAPWR.n44 VAPWR.t38 707.519
R39 VAPWR.n47 VAPWR.t36 707.519
R40 VAPWR.n4 VAPWR.t24 707.519
R41 VAPWR.n2 VAPWR.t40 707.519
R42 VAPWR.n61 VAPWR.n60 13.3797
R43 VAPWR.n58 VAPWR.n57 13.3797
R44 VAPWR.n33 VAPWR.n32 13.3797
R45 VAPWR.n8 VAPWR.n7 13.3797
R46 VAPWR.n12 VAPWR.n11 13.3797
R47 VAPWR.n23 VAPWR.n22 13.3797
R48 VAPWR.n20 VAPWR.n19 13.3797
R49 VAPWR.n17 VAPWR.n16 13.3797
R50 VAPWR.n14 VAPWR.n13 13.3797
R51 VAPWR.n10 VAPWR.n9 13.3797
R52 VAPWR.n28 VAPWR.n27 13.3797
R53 VAPWR.n53 VAPWR.n52 13.3223
R54 VAPWR VAPWR.n54 13.3223
R55 VAPWR.n39 VAPWR.n38 13.3223
R56 VAPWR.n35 VAPWR.n34 13.3223
R57 VAPWR VAPWR.n6 13.3223
R58 VAPWR.n42 VAPWR.n41 13.3223
R59 VAPWR.n45 VAPWR.n44 13.3223
R60 VAPWR.n48 VAPWR.n47 13.3223
R61 VAPWR.n5 VAPWR.n4 13.3223
R62 VAPWR.n3 VAPWR.n2 13.3223
R63 VAPWR.n59 VAPWR.n58 9.70762
R64 VAPWR.n18 VAPWR.n15 9.45042
R65 VAPWR.n31 VAPWR 8.52916
R66 VAPWR.n62 VAPWR.n61 7.92611
R67 VAPWR.n40 VAPWR.n37 7.71912
R68 VAPWR.n15 VAPWR.n14 7.71771
R69 VAPWR.n31 VAPWR.n30 7.41572
R70 VAPWR.n55 VAPWR 7.13154
R71 VAPWR.n40 VAPWR.n39 7.11663
R72 VAPWR.n18 VAPWR.n17 7.10884
R73 VAPWR.n43 VAPWR.n42 6.89753
R74 VAPWR.n21 VAPWR.n20 6.54898
R75 VAPWR.n49 VAPWR.n46 6.23852
R76 VAPWR.n30 VAPWR.n8 6.19396
R77 VAPWR.n46 VAPWR.n45 6.10554
R78 VAPWR.n29 VAPWR.n28 6.01845
R79 VAPWR.n36 VAPWR.n35 5.92055
R80 VAPWR.n49 VAPWR.n48 5.84717
R81 VAPWR.n24 VAPWR.n23 5.78073
R82 VAPWR.n26 VAPWR.n10 5.73072
R83 VAPWR.n50 VAPWR.n5 5.60146
R84 VAPWR.n51 VAPWR.n3 5.59565
R85 VAPWR.n25 VAPWR.n12 5.50466
R86 VAPWR.n55 VAPWR.n53 4.89777
R87 VAPWR.n36 VAPWR.n33 4.86074
R88 VAPWR.n46 VAPWR.n43 4.01511
R89 VAPWR.n66 VAPWR 3.49767
R90 VAPWR.n67 VAPWR 3.44936
R91 VAPWR.n37 VAPWR.n36 2.91269
R92 VAPWR.n59 VAPWR.n56 2.82184
R93 VAPWR.n1 VAPWR.n0 1.63622
R94 VAPWR.n24 VAPWR.n21 1.36014
R95 VAPWR.n30 VAPWR.n29 1.34127
R96 VAPWR.n56 VAPWR.n51 1.32921
R97 VAPWR.n56 VAPWR.n55 1.313
R98 VAPWR.n63 VAPWR.n0 1.29727
R99 VAPWR.n29 VAPWR.n26 1.10191
R100 VAPWR.n51 VAPWR.n50 0.940035
R101 VAPWR.n62 VAPWR.n59 0.85748
R102 VAPWR.n37 VAPWR.n31 0.767594
R103 VAPWR.n66 VAPWR.n65 0.616014
R104 VAPWR.n25 VAPWR.n24 0.52495
R105 VAPWR.n43 VAPWR.n40 0.514977
R106 VAPWR.n15 VAPWR.n1 0.507476
R107 VAPWR.n26 VAPWR.n25 0.505442
R108 VAPWR.n21 VAPWR.n18 0.500622
R109 VAPWR.n50 VAPWR.n49 0.483622
R110 VAPWR.n65 VAPWR.n0 0.20333
R111 VAPWR VAPWR.n67 0.193138
R112 VAPWR.n61 VAPWR 0.057877
R113 VAPWR.n58 VAPWR 0.057877
R114 VAPWR.n33 VAPWR 0.057877
R115 VAPWR.n8 VAPWR 0.057877
R116 VAPWR.n12 VAPWR 0.057877
R117 VAPWR.n23 VAPWR 0.057877
R118 VAPWR.n20 VAPWR 0.057877
R119 VAPWR.n17 VAPWR 0.057877
R120 VAPWR.n14 VAPWR 0.057877
R121 VAPWR.n10 VAPWR 0.057877
R122 VAPWR.n28 VAPWR 0.057877
R123 VAPWR.n53 VAPWR 0.0496071
R124 VAPWR.n39 VAPWR 0.0496071
R125 VAPWR.n35 VAPWR 0.0496071
R126 VAPWR.n42 VAPWR 0.0496071
R127 VAPWR.n45 VAPWR 0.0496071
R128 VAPWR.n48 VAPWR 0.0496071
R129 VAPWR.n5 VAPWR 0.0496071
R130 VAPWR.n3 VAPWR 0.0496071
R131 VAPWR.n65 VAPWR.n64 0.0335189
R132 VAPWR.n64 VAPWR.n1 0.00474612
R133 VAPWR.n63 VAPWR.n62 0.00305102
R134 VAPWR.n64 VAPWR.n63 0.00285849
R135 VAPWR.n67 VAPWR.n66 0.0018126
R136 VGND.n194 VGND.n193 101372
R137 VGND.n141 VGND.n140 97829.8
R138 VGND.n452 VGND.n9 64989.2
R139 VGND.n232 VGND.n144 63317.7
R140 VGND.n196 VGND.n173 51969.6
R141 VGND.n286 VGND.n285 50528.4
R142 VGND.n238 VGND.n145 49981.2
R143 VGND.n236 VGND.t0 48989.1
R144 VGND.n195 VGND.n153 48956.8
R145 VGND.n116 VGND.n14 46397.1
R146 VGND.n242 VGND.n240 34056.2
R147 VGND.n285 VGND.t61 32820.9
R148 VGND.n201 VGND.n196 31013.9
R149 VGND.n410 VGND.n26 29705.2
R150 VGND.n238 VGND.n146 26125.9
R151 VGND.n236 VGND.n235 24501.8
R152 VGND.n233 VGND.n146 22668.4
R153 VGND.n195 VGND.n194 20954.6
R154 VGND.n140 VGND.n26 20954.6
R155 VGND.n237 VGND.n12 18294.4
R156 VGND.t84 VGND.n14 14642.2
R157 VGND.n196 VGND.n195 13862.9
R158 VGND.n285 VGND.n26 13853.3
R159 VGND.n181 VGND.n177 12938.5
R160 VGND.n236 VGND.n146 10983.3
R161 VGND.n116 VGND.n115 10461.7
R162 VGND.n232 VGND.t48 8761.83
R163 VGND.n234 VGND.n233 8254.98
R164 VGND.n175 VGND.n173 8219.71
R165 VGND.n140 VGND.n9 8171.07
R166 VGND.n194 VGND.n144 8164.43
R167 VGND.n453 VGND.n452 8158.04
R168 VGND.n452 VGND.n12 8007.21
R169 VGND.n233 VGND.n232 8000.6
R170 VGND.n143 VGND.n139 7798.05
R171 VGND.n116 VGND 7183.82
R172 VGND.n238 VGND.n144 6658.85
R173 VGND.n12 VGND.n11 6298.11
R174 VGND.n180 VGND.n177 5767.96
R175 VGND.n232 VGND.n153 5608.83
R176 VGND.n284 VGND.n141 5496.81
R177 VGND.n409 VGND.n408 5446.6
R178 VGND.n182 VGND.n181 5163.17
R179 VGND.n240 VGND.n9 4690.48
R180 VGND.n235 VGND.n147 4323.23
R181 VGND.n150 VGND.n12 4311.21
R182 VGND.n286 VGND.n284 4138.55
R183 VGND.n193 VGND.n192 3936.62
R184 VGND.n241 VGND.n141 3888.93
R185 VGND.n192 VGND.n145 3732.38
R186 VGND.n190 VGND.n177 3431.95
R187 VGND.n181 VGND.n143 3199.08
R188 VGND.n239 VGND.n143 3097.77
R189 VGND.n238 VGND.n237 3097.77
R190 VGND.n191 VGND.n176 3043.22
R191 VGND.n180 VGND.n179 3033.4
R192 VGND.t80 VGND.n139 2956.47
R193 VGND.n242 VGND.n241 2771.85
R194 VGND.n152 VGND.n150 2374.28
R195 VGND.n150 VGND.n149 2325.64
R196 VGND.n193 VGND.t23 2293.69
R197 VGND.n452 VGND.n13 2139.51
R198 VGND.t48 VGND.n231 2108.34
R199 VGND.n191 VGND.n143 2021.45
R200 VGND.t7 VGND.n180 1675.99
R201 VGND.n11 VGND.t2 1523.34
R202 VGND.n453 VGND.t11 1523.34
R203 VGND.n176 VGND.t52 1523.34
R204 VGND.n286 VGND.n139 1501.79
R205 VGND.n191 VGND.n173 1498.22
R206 VGND.n141 VGND.t76 1467.82
R207 VGND.n193 VGND.n175 1415.65
R208 VGND.t96 VGND.n153 1206.01
R209 VGND.n414 VGND.n413 1198.25
R210 VGND.n412 VGND.n24 1198.25
R211 VGND.n242 VGND.t80 1186.75
R212 VGND.n192 VGND.n191 1105.93
R213 VGND.n292 VGND.t32 958.28
R214 VGND.n243 VGND.n242 921.593
R215 VGND.n182 VGND.t7 912.855
R216 VGND.t88 VGND.n203 905.449
R217 VGND.t59 VGND.n198 842.21
R218 VGND.t92 VGND.t63 809.293
R219 VGND.t94 VGND.t90 800.774
R220 VGND.n241 VGND.n139 754.139
R221 VGND.n451 VGND.n14 613.852
R222 VGND.n115 VGND.n114 595.942
R223 VGND.t65 VGND.n286 592.851
R224 VGND.n198 VGND.n197 585
R225 VGND.n200 VGND.n199 585
R226 VGND.n451 VGND.n450 585
R227 VGND.n11 VGND.n10 585
R228 VGND.n149 VGND.n148 585
R229 VGND.n152 VGND.n151 585
R230 VGND.n454 VGND.n453 585
R231 VGND.n335 VGND.n13 585
R232 VGND.n293 VGND.n292 585
R233 VGND.n291 VGND.n290 585
R234 VGND.n408 VGND.n407 585
R235 VGND.n284 VGND.n283 585
R236 VGND.n175 VGND.n174 585
R237 VGND.n203 VGND.n202 585
R238 VGND.n205 VGND.n204 585
R239 VGND.n186 VGND.n176 585
R240 VGND.n190 VGND.n189 585
R241 VGND.n183 VGND.n182 585
R242 VGND.n179 VGND.n178 585
R243 VGND.n149 VGND.t0 574.539
R244 VGND.t86 VGND.n201 533.332
R245 VGND.n408 VGND.t61 489.839
R246 VGND.n204 VGND.n173 489.707
R247 VGND.t36 VGND.t72 451.5
R248 VGND.t38 VGND.t36 430.204
R249 VGND.t82 VGND.n234 424.175
R250 VGND.t72 VGND.t92 404.647
R251 VGND.t90 VGND.t84 404.647
R252 VGND.n201 VGND.n200 382.728
R253 VGND.n411 VGND.t38 370.572
R254 VGND.t15 VGND.n152 362.452
R255 VGND.t52 VGND.n145 360.884
R256 VGND.t63 VGND.t94 357.793
R257 VGND.n452 VGND.t13 313.435
R258 VGND.n183 VGND.t8 282.13
R259 VGND.n243 VGND.t81 282.13
R260 VGND.n407 VGND.t62 282.13
R261 VGND.n148 VGND.t1 282.13
R262 VGND.n10 VGND.t3 282.13
R263 VGND.n151 VGND.t16 282.13
R264 VGND.n454 VGND.t12 282.13
R265 VGND.n335 VGND.t27 282.13
R266 VGND.n290 VGND.t33 282.13
R267 VGND.n293 VGND.t66 282.13
R268 VGND.n283 VGND.t77 282.13
R269 VGND.n450 VGND.t14 281.841
R270 VGND.n231 VGND.t49 281.839
R271 VGND.n199 VGND.t60 281.839
R272 VGND.n197 VGND.t97 281.839
R273 VGND.n186 VGND.t53 281.839
R274 VGND.n189 VGND.t51 281.839
R275 VGND.n147 VGND.t83 281.839
R276 VGND.n178 VGND.t21 281.839
R277 VGND.n174 VGND.t24 281.839
R278 VGND.n205 VGND.t89 281.839
R279 VGND.n202 VGND.t87 281.839
R280 VGND.n237 VGND.n236 264.286
R281 VGND.n90 VGND.t45 251
R282 VGND.n57 VGND.t68 251
R283 VGND.n437 VGND.t93 251
R284 VGND.n234 VGND.t15 245.631
R285 VGND.n104 VGND.t25 243.028
R286 VGND.n44 VGND.t58 243.028
R287 VGND.n424 VGND.t79 243.028
R288 VGND.n411 VGND.t26 232.994
R289 VGND.n77 VGND.n76 218.506
R290 VGND.n59 VGND.n58 218.506
R291 VGND.n439 VGND.n438 218.506
R292 VGND.t13 VGND.n451 212.357
R293 VGND.n239 VGND.n238 209.014
R294 VGND.n80 VGND.n79 200.201
R295 VGND.n66 VGND.n30 200.201
R296 VGND.n447 VGND.n446 200.201
R297 VGND.n108 VGND.n70 199.739
R298 VGND.n40 VGND.n39 199.739
R299 VGND.n420 VGND.n419 199.739
R300 VGND.n98 VGND.n97 199.53
R301 VGND.n50 VGND.n35 199.53
R302 VGND.n430 VGND.n21 199.53
R303 VGND.t26 VGND.n13 196.702
R304 VGND.n409 VGND.n116 165.179
R305 VGND.n292 VGND.t65 162.868
R306 VGND.t32 VGND.n291 162.868
R307 VGND.n204 VGND.t88 153.888
R308 VGND.n203 VGND.t86 153.888
R309 VGND.n200 VGND.t59 151.095
R310 VGND.n198 VGND.t96 151.095
R311 VGND.n191 VGND.t50 130.082
R312 VGND.t20 VGND.n139 129.425
R313 VGND.t6 VGND 118.189
R314 VGND.t50 VGND.n190 99.8351
R315 VGND.n179 VGND.t20 99.332
R316 VGND.n97 VGND.t37 74.8666
R317 VGND.n35 VGND.t5 74.8666
R318 VGND.n21 VGND.t39 74.8666
R319 VGND.t28 VGND.t44 69.615
R320 VGND.t40 VGND.t42 68.8822
R321 VGND.t74 VGND.t78 68.8822
R322 VGND.n235 VGND.t82 54.4208
R323 VGND.n79 VGND.t41 54.2862
R324 VGND.n30 VGND.t67 54.2862
R325 VGND.n446 VGND.t91 54.2862
R326 VGND.n291 VGND.n116 53.7948
R327 VGND.t78 VGND.t73 41.0364
R328 VGND.n97 VGND.t17 40.0005
R329 VGND.n35 VGND.t10 40.0005
R330 VGND.n21 VGND.t71 40.0005
R331 VGND.t46 VGND.t34 38.838
R332 VGND.n70 VGND.t22 38.5719
R333 VGND.n70 VGND.t47 38.5719
R334 VGND.n39 VGND.t31 38.5719
R335 VGND.n39 VGND.t30 38.5719
R336 VGND.n419 VGND.t19 38.5719
R337 VGND.n419 VGND.t75 38.5719
R338 VGND.t73 VGND.t35 36.2733
R339 VGND.t35 VGND.t70 36.2733
R340 VGND.t44 VGND.t46 34.8077
R341 VGND.t54 VGND.t40 34.8077
R342 VGND.n86 VGND.n85 34.6358
R343 VGND.n85 VGND.n84 34.6358
R344 VGND.n96 VGND.n95 34.6358
R345 VGND.n95 VGND.n74 34.6358
R346 VGND.n91 VGND.n74 34.6358
R347 VGND.n103 VGND.n102 34.6358
R348 VGND.n102 VGND.n72 34.6358
R349 VGND.n64 VGND.n31 34.6358
R350 VGND.n65 VGND.n64 34.6358
R351 VGND.n52 VGND.n51 34.6358
R352 VGND.n52 VGND.n33 34.6358
R353 VGND.n56 VGND.n33 34.6358
R354 VGND.n45 VGND.n37 34.6358
R355 VGND.n49 VGND.n37 34.6358
R356 VGND.n426 VGND.n425 34.6358
R357 VGND.n426 VGND.n20 34.6358
R358 VGND.n432 VGND.n431 34.6358
R359 VGND.n432 VGND.n18 34.6358
R360 VGND.n436 VGND.n18 34.6358
R361 VGND.n444 VGND.n16 34.6358
R362 VGND.n445 VGND.n444 34.6358
R363 VGND.n413 VGND.n412 33.7085
R364 VGND.n412 VGND 33.7085
R365 VGND.n89 VGND.n77 32.7534
R366 VGND.n60 VGND.n59 32.7534
R367 VGND.n440 VGND.n439 32.7534
R368 VGND.t4 VGND.t9 31.3274
R369 VGND.n90 VGND.n89 31.2476
R370 VGND.n60 VGND.n57 31.2476
R371 VGND.n440 VGND.n437 31.2476
R372 VGND.n98 VGND.n72 30.8711
R373 VGND.n50 VGND.n49 30.8711
R374 VGND.n430 VGND.n20 30.8711
R375 VGND.t42 VGND.t28 30.7774
R376 VGND.t18 VGND.t74 30.7774
R377 VGND.n104 VGND.n103 27.4829
R378 VGND.n45 VGND.n44 27.4829
R379 VGND.n425 VGND.n424 27.4829
R380 VGND.n79 VGND.t55 25.9346
R381 VGND.n30 VGND.t98 25.9346
R382 VGND.n446 VGND.t85 25.9346
R383 VGND.n410 VGND.t54 25.6479
R384 VGND.n413 VGND.n410 25.6479
R385 VGND.n76 VGND.t29 24.9236
R386 VGND.n76 VGND.t43 24.9236
R387 VGND.n58 VGND.t57 24.9236
R388 VGND.n58 VGND.t69 24.9236
R389 VGND.n438 VGND.t64 24.9236
R390 VGND.n438 VGND.t95 24.9236
R391 VGND.n187 VGND.n172 23.8791
R392 VGND.n414 VGND.n25 23.7181
R393 VGND.n84 VGND.n80 23.7181
R394 VGND.n109 VGND.n27 23.7181
R395 VGND.n113 VGND.n28 23.7181
R396 VGND.n66 VGND.n65 23.7181
R397 VGND.n418 VGND.n24 23.7181
R398 VGND.n447 VGND.n445 23.7181
R399 VGND.n230 VGND.n1 23.1262
R400 VGND.n108 VGND.n69 22.9652
R401 VGND.n104 VGND.n69 22.9652
R402 VGND.n43 VGND.n40 22.9652
R403 VGND.n44 VGND.n43 22.9652
R404 VGND.n420 VGND.n23 22.9652
R405 VGND.n424 VGND.n23 22.9652
R406 VGND.n115 VGND.t56 22.7837
R407 VGND.n91 VGND.n90 22.2123
R408 VGND.n57 VGND.n56 22.2123
R409 VGND.n437 VGND.n436 22.2123
R410 VGND.n80 VGND.n25 21.4593
R411 VGND.n109 VGND.n108 21.4593
R412 VGND.n66 VGND.n28 21.4593
R413 VGND.n420 VGND.n418 21.4593
R414 VGND.n462 VGND.n461 20.8917
R415 VGND.n245 VGND.n142 19.445
R416 VGND.n240 VGND.n239 15.7795
R417 VGND.n184 VGND.n183 13.2958
R418 VGND.n244 VGND.n243 13.2958
R419 VGND.n407 VGND.n406 13.2958
R420 VGND.n148 VGND.n3 13.2958
R421 VGND.n10 VGND.n4 13.2958
R422 VGND.n151 VGND.n2 13.2958
R423 VGND.n455 VGND.n454 13.2958
R424 VGND.n336 VGND.n335 13.2958
R425 VGND.n290 VGND.n289 13.2958
R426 VGND.n294 VGND.n293 13.2958
R427 VGND.n283 VGND.n282 13.2958
R428 VGND.n197 VGND 13.2396
R429 VGND.n199 VGND 13.2396
R430 VGND VGND.n186 13.2396
R431 VGND.n189 VGND 13.2396
R432 VGND.n450 VGND 13.2396
R433 VGND.n147 VGND 13.2396
R434 VGND.n178 VGND 13.2396
R435 VGND.n174 VGND 13.2396
R436 VGND VGND.n205 13.2396
R437 VGND.n202 VGND 13.2396
R438 VGND.n231 VGND 13.2396
R439 VGND.t34 VGND.n409 13.1906
R440 VGND VGND.n449 12.8296
R441 VGND.n414 VGND.n24 12.8005
R442 VGND.n449 VGND 12.1807
R443 VGND.t70 VGND.n411 11.725
R444 VGND.n188 VGND.n187 11.3685
R445 VGND VGND.t18 11.3586
R446 VGND.n98 VGND.n96 10.5417
R447 VGND.n51 VGND.n50 10.5417
R448 VGND.n431 VGND.n430 10.5417
R449 VGND.n445 VGND.n15 9.3005
R450 VGND.n444 VGND.n443 9.3005
R451 VGND.n442 VGND.n16 9.3005
R452 VGND.n441 VGND.n440 9.3005
R453 VGND.n437 VGND.n17 9.3005
R454 VGND.n436 VGND.n435 9.3005
R455 VGND.n434 VGND.n18 9.3005
R456 VGND.n433 VGND.n432 9.3005
R457 VGND.n431 VGND.n19 9.3005
R458 VGND.n430 VGND.n429 9.3005
R459 VGND.n428 VGND.n20 9.3005
R460 VGND.n427 VGND.n426 9.3005
R461 VGND.n425 VGND.n22 9.3005
R462 VGND.n424 VGND.n423 9.3005
R463 VGND.n422 VGND.n23 9.3005
R464 VGND.n421 VGND.n420 9.3005
R465 VGND.n418 VGND.n417 9.3005
R466 VGND.n416 VGND.n24 9.3005
R467 VGND.n43 VGND.n42 9.3005
R468 VGND.n44 VGND.n38 9.3005
R469 VGND.n46 VGND.n45 9.3005
R470 VGND.n47 VGND.n37 9.3005
R471 VGND.n49 VGND.n48 9.3005
R472 VGND.n50 VGND.n36 9.3005
R473 VGND.n51 VGND.n34 9.3005
R474 VGND.n53 VGND.n52 9.3005
R475 VGND.n54 VGND.n33 9.3005
R476 VGND.n56 VGND.n55 9.3005
R477 VGND.n57 VGND.n32 9.3005
R478 VGND.n61 VGND.n60 9.3005
R479 VGND.n62 VGND.n31 9.3005
R480 VGND.n64 VGND.n63 9.3005
R481 VGND.n65 VGND.n29 9.3005
R482 VGND.n67 VGND.n66 9.3005
R483 VGND.n68 VGND.n28 9.3005
R484 VGND.n113 VGND.n112 9.3005
R485 VGND.n111 VGND.n27 9.3005
R486 VGND.n110 VGND.n109 9.3005
R487 VGND.n108 VGND.n107 9.3005
R488 VGND.n106 VGND.n69 9.3005
R489 VGND.n105 VGND.n104 9.3005
R490 VGND.n103 VGND.n71 9.3005
R491 VGND.n102 VGND.n101 9.3005
R492 VGND.n100 VGND.n72 9.3005
R493 VGND.n99 VGND.n98 9.3005
R494 VGND.n96 VGND.n73 9.3005
R495 VGND.n95 VGND.n94 9.3005
R496 VGND.n93 VGND.n74 9.3005
R497 VGND.n92 VGND.n91 9.3005
R498 VGND.n90 VGND.n75 9.3005
R499 VGND.n89 VGND.n88 9.3005
R500 VGND.n87 VGND.n86 9.3005
R501 VGND.n85 VGND.n78 9.3005
R502 VGND.n84 VGND.n83 9.3005
R503 VGND.n82 VGND.n80 9.3005
R504 VGND.n81 VGND.n25 9.3005
R505 VGND.n415 VGND.n414 9.3005
R506 VGND VGND.n1 9.06372
R507 VGND.t9 VGND.t6 8.54419
R508 VGND.n185 VGND.n184 7.79935
R509 VGND.n245 VGND.n244 7.42221
R510 VGND.n41 VGND.n40 7.12576
R511 VGND.n448 VGND.n447 7.12063
R512 VGND.n463 VGND.n3 6.96
R513 VGND VGND.n230 6.82321
R514 VGND.n114 VGND.n113 6.367
R515 VGND.n114 VGND.n27 6.367
R516 VGND.n464 VGND.n2 6.32363
R517 VGND.n282 VGND.n281 6.24462
R518 VGND.n228 VGND 6.10287
R519 VGND VGND.n142 5.99098
R520 VGND.n187 VGND 5.98182
R521 VGND.n462 VGND.n4 5.94997
R522 VGND.n456 VGND.n455 5.91022
R523 VGND VGND.n172 5.81859
R524 VGND.n289 VGND.n288 5.80858
R525 VGND.n295 VGND.n294 5.70662
R526 VGND VGND.n171 5.69376
R527 VGND.n206 VGND 5.57954
R528 VGND.n207 VGND 5.53239
R529 VGND VGND.n188 5.49935
R530 VGND.n382 VGND.n336 5.39911
R531 VGND.n119 VGND.n118 5.04217
R532 VGND.n406 VGND.n405 5.00883
R533 VGND.n449 VGND.n0 4.99159
R534 VGND.n0 VGND 3.44325
R535 VGND.n467 VGND 3.36335
R536 VGND.n316 VGND.n118 3.29217
R537 VGND.n246 VGND.n245 3.10947
R538 VGND VGND.n467 2.3855
R539 VGND.n86 VGND.n77 1.88285
R540 VGND.n59 VGND.n31 1.88285
R541 VGND.n439 VGND.n16 1.88285
R542 VGND.n372 VGND.n371 1.5618
R543 VGND.t56 VGND.t4 1.42445
R544 VGND.n405 VGND.n117 1.2755
R545 VGND.n188 VGND.n185 1.26584
R546 VGND.n288 VGND.n287 0.979021
R547 VGND.n230 VGND.n229 0.96878
R548 VGND.n464 VGND.n463 0.964749
R549 VGND.n185 VGND.n142 0.956896
R550 VGND.n463 VGND.n462 0.903134
R551 VGND.n207 VGND.n206 0.844578
R552 VGND.n371 VGND.n370 0.777168
R553 VGND.n466 VGND.n465 0.726602
R554 VGND.n206 VGND.n172 0.707232
R555 VGND.n288 VGND.n118 0.6755
R556 VGND.n405 VGND.n404 0.638
R557 VGND.n208 VGND.n207 0.577069
R558 VGND.n287 VGND.n120 0.574766
R559 VGND.n465 VGND.n1 0.561048
R560 VGND.n370 VGND.n369 0.533644
R561 VGND.n121 VGND.n120 0.469554
R562 VGND.n122 VGND.n121 0.431514
R563 VGND.n317 VGND.n316 0.425271
R564 VGND.n369 VGND.n368 0.420347
R565 VGND.n368 VGND.n367 0.36938
R566 VGND.n123 VGND.n122 0.355217
R567 VGND.n367 VGND.n366 0.332442
R568 VGND.n124 VGND.n123 0.314827
R569 VGND.n209 VGND.n208 0.307815
R570 VGND.n366 VGND.n365 0.293921
R571 VGND.n125 VGND.n124 0.283145
R572 VGND.n365 VGND.n364 0.262603
R573 VGND.n126 VGND.n125 0.257575
R574 VGND.n364 VGND.n363 0.242676
R575 VGND.n127 VGND.n126 0.242107
R576 VGND.n363 VGND.n362 0.227688
R577 VGND.n128 VGND.n127 0.224203
R578 VGND.n295 VGND.n138 0.21925
R579 VGND.n362 VGND.n361 0.214493
R580 VGND.n129 VGND.n128 0.209128
R581 VGND.n229 VGND.n154 0.207265
R582 VGND.n361 VGND.n357 0.207112
R583 VGND.n362 VGND.n356 0.205418
R584 VGND.n363 VGND.n355 0.203752
R585 VGND.n210 VGND.n209 0.202174
R586 VGND.n361 VGND.n360 0.201991
R587 VGND.n364 VGND.n354 0.2005
R588 VGND.n365 VGND.n353 0.198913
R589 VGND.n366 VGND.n352 0.19735
R590 VGND.n130 VGND.n129 0.196195
R591 VGND.n367 VGND.n351 0.195812
R592 VGND.n360 VGND.n8 0.194723
R593 VGND.n368 VGND.n350 0.194298
R594 VGND.n456 VGND.n7 0.193682
R595 VGND.n369 VGND.n349 0.19134
R596 VGND.n211 VGND.n210 0.190823
R597 VGND.n370 VGND.n348 0.189894
R598 VGND.n131 VGND.n130 0.189066
R599 VGND.n371 VGND.n347 0.18847
R600 VGND.n461 VGND.n5 0.188059
R601 VGND.n212 VGND.n211 0.184664
R602 VGND.n460 VGND.n459 0.181056
R603 VGND.n213 VGND.n212 0.180457
R604 VGND.n132 VGND.n131 0.179109
R605 VGND.n133 VGND.n132 0.178762
R606 VGND.n214 VGND.n213 0.167949
R607 VGND.n134 VGND.n133 0.166149
R608 VGND.n281 VGND.n246 0.165057
R609 VGND.n216 VGND.n215 0.164532
R610 VGND.n215 VGND.n214 0.164276
R611 VGND.n136 VGND.n135 0.159573
R612 VGND.n400 VGND.n399 0.159247
R613 VGND.n135 VGND.n134 0.159247
R614 VGND.n381 VGND.n380 0.156646
R615 VGND.n399 VGND.n398 0.156448
R616 VGND.n217 VGND.n216 0.155102
R617 VGND.n314 VGND.n120 0.154588
R618 VGND.n360 VGND.n359 0.153861
R619 VGND.n313 VGND.n121 0.153802
R620 VGND.n296 VGND.n136 0.153257
R621 VGND.n218 VGND.n217 0.153062
R622 VGND.n312 VGND.n122 0.153016
R623 VGND VGND.n448 0.152603
R624 VGND.n400 VGND.n117 0.152527
R625 VGND.n310 VGND.n124 0.152399
R626 VGND.n404 VGND.n317 0.152332
R627 VGND.n311 VGND.n123 0.15223
R628 VGND.n397 VGND.n396 0.151068
R629 VGND.n308 VGND.n126 0.150816
R630 VGND.n219 VGND.n218 0.150802
R631 VGND.n309 VGND.n125 0.150657
R632 VGND.n398 VGND.n397 0.15035
R633 VGND.n306 VGND.n128 0.150182
R634 VGND.n226 VGND.n225 0.150148
R635 VGND.n307 VGND.n127 0.150025
R636 VGND.n209 VGND.n170 0.149538
R637 VGND.n305 VGND.n129 0.149385
R638 VGND.n211 VGND.n168 0.148887
R639 VGND.n210 VGND.n169 0.148737
R640 VGND.n304 VGND.n130 0.148589
R641 VGND.n448 VGND.n15 0.148519
R642 VGND.n212 VGND.n167 0.148081
R643 VGND.n302 VGND.n132 0.147936
R644 VGND.n303 VGND.n131 0.147793
R645 VGND.n215 VGND.n164 0.147559
R646 VGND.n315 VGND.n119 0.147513
R647 VGND.n214 VGND.n165 0.147416
R648 VGND.n401 VGND.n400 0.147274
R649 VGND.n300 VGND.n134 0.147274
R650 VGND.n213 VGND.n166 0.147274
R651 VGND.n403 VGND.n402 0.147135
R652 VGND.n301 VGND.n133 0.147135
R653 VGND.n218 VGND.n161 0.147023
R654 VGND.n373 VGND.n345 0.146955
R655 VGND.n216 VGND.n163 0.146742
R656 VGND.n399 VGND.n318 0.146468
R657 VGND.n299 VGND.n135 0.146468
R658 VGND.n219 VGND.n160 0.146195
R659 VGND.n220 VGND.n219 0.146195
R660 VGND.n396 VGND.n395 0.146191
R661 VGND.n262 VGND.n138 0.146191
R662 VGND.n396 VGND.n321 0.145925
R663 VGND.n138 VGND.n137 0.145925
R664 VGND.n217 VGND.n162 0.145925
R665 VGND.n397 VGND.n320 0.145792
R666 VGND.n297 VGND.n296 0.145792
R667 VGND.n223 VGND.n156 0.14577
R668 VGND.n224 VGND.n155 0.14577
R669 VGND.n398 VGND.n319 0.145661
R670 VGND.n298 VGND.n136 0.145661
R671 VGND.n222 VGND.n157 0.145634
R672 VGND.n375 VGND.n343 0.145573
R673 VGND.n221 VGND.n158 0.1455
R674 VGND.n376 VGND.n342 0.145428
R675 VGND.n393 VGND.n324 0.145368
R676 VGND.n264 VGND.n259 0.145368
R677 VGND.n220 VGND.n159 0.145368
R678 VGND.n377 VGND.n341 0.145284
R679 VGND.n395 VGND.n322 0.145108
R680 VGND.n262 VGND.n261 0.145108
R681 VGND.n277 VGND.n276 0.144866
R682 VGND.n389 VGND.n328 0.144795
R683 VGND.n268 VGND.n255 0.144795
R684 VGND.n221 VGND.n220 0.144667
R685 VGND.n374 VGND.n344 0.144661
R686 VGND.n392 VGND.n325 0.14454
R687 VGND.n265 VGND.n258 0.14454
R688 VGND.n273 VGND.n250 0.144466
R689 VGND.n385 VGND.n332 0.144336
R690 VGND.n272 VGND.n251 0.144336
R691 VGND.n394 VGND.n323 0.144291
R692 VGND.n263 VGND.n260 0.144291
R693 VGND.n378 VGND.n340 0.14425
R694 VGND.n379 VGND.n339 0.144117
R695 VGND.n280 VGND.n279 0.144117
R696 VGND.n387 VGND.n330 0.144081
R697 VGND.n388 VGND.n329 0.144081
R698 VGND.n270 VGND.n253 0.144081
R699 VGND.n269 VGND.n254 0.144081
R700 VGND.n380 VGND.n338 0.143986
R701 VGND.n278 VGND.n247 0.143986
R702 VGND.n390 VGND.n327 0.143833
R703 VGND.n267 VGND.n256 0.143833
R704 VGND.n275 VGND.n248 0.143729
R705 VGND.n391 VGND.n326 0.143712
R706 VGND.n266 VGND.n257 0.143712
R707 VGND.n274 VGND.n249 0.143603
R708 VGND.n42 VGND.n41 0.143396
R709 VGND.n386 VGND.n331 0.143357
R710 VGND.n271 VGND.n252 0.143357
R711 VGND.n222 VGND.n221 0.143343
R712 VGND.n394 VGND.n393 0.142608
R713 VGND.n264 VGND.n263 0.142608
R714 VGND.n223 VGND.n222 0.142204
R715 VGND.n395 VGND.n394 0.14174
R716 VGND.n263 VGND.n262 0.14174
R717 VGND.n227 VGND.n154 0.141228
R718 VGND.n225 VGND.n224 0.140944
R719 VGND.n224 VGND.n223 0.14022
R720 VGND.n225 VGND.n154 0.139918
R721 VGND.n393 VGND.n392 0.138984
R722 VGND.n265 VGND.n264 0.138984
R723 VGND.n268 VGND.n267 0.137868
R724 VGND.n266 VGND.n265 0.137764
R725 VGND.n267 VGND.n266 0.13669
R726 VGND.n390 VGND.n389 0.135675
R727 VGND.n392 VGND.n391 0.135449
R728 VGND.n374 VGND.n373 0.134751
R729 VGND.n391 VGND.n390 0.134458
R730 VGND.n270 VGND.n269 0.134444
R731 VGND.n272 VGND.n271 0.13348
R732 VGND.n375 VGND.n374 0.133147
R733 VGND.n388 VGND.n387 0.132395
R734 VGND.n389 VGND.n388 0.132323
R735 VGND.n269 VGND.n268 0.132323
R736 VGND.n274 VGND.n273 0.131889
R737 VGND.n276 VGND.n247 0.131852
R738 VGND.n378 VGND.n377 0.13184
R739 VGND.n280 VGND.n247 0.131755
R740 VGND.n376 VGND.n375 0.131611
R741 VGND.n276 VGND.n275 0.131576
R742 VGND.n386 VGND.n385 0.131557
R743 VGND.n271 VGND.n270 0.131307
R744 VGND.n377 VGND.n376 0.131251
R745 VGND.n385 VGND.n384 0.130509
R746 VGND.n273 VGND.n272 0.130509
R747 VGND.n379 VGND.n378 0.130342
R748 VGND.n275 VGND.n274 0.130162
R749 VGND.n380 VGND.n379 0.13011
R750 VGND.n384 VGND.n383 0.130051
R751 VGND.n387 VGND.n386 0.129353
R752 VGND.n346 VGND.n345 0.124567
R753 VGND.n42 VGND.n38 0.120292
R754 VGND.n46 VGND.n38 0.120292
R755 VGND.n47 VGND.n46 0.120292
R756 VGND.n48 VGND.n47 0.120292
R757 VGND.n48 VGND.n36 0.120292
R758 VGND.n36 VGND.n34 0.120292
R759 VGND.n53 VGND.n34 0.120292
R760 VGND.n54 VGND.n53 0.120292
R761 VGND.n55 VGND.n54 0.120292
R762 VGND.n55 VGND.n32 0.120292
R763 VGND.n61 VGND.n32 0.120292
R764 VGND.n62 VGND.n61 0.120292
R765 VGND.n63 VGND.n62 0.120292
R766 VGND.n63 VGND.n29 0.120292
R767 VGND.n67 VGND.n29 0.120292
R768 VGND.n68 VGND.n67 0.120292
R769 VGND.n107 VGND.n106 0.120292
R770 VGND.n106 VGND.n105 0.120292
R771 VGND.n105 VGND.n71 0.120292
R772 VGND.n101 VGND.n71 0.120292
R773 VGND.n101 VGND.n100 0.120292
R774 VGND.n100 VGND.n99 0.120292
R775 VGND.n99 VGND.n73 0.120292
R776 VGND.n94 VGND.n73 0.120292
R777 VGND.n94 VGND.n93 0.120292
R778 VGND.n93 VGND.n92 0.120292
R779 VGND.n92 VGND.n75 0.120292
R780 VGND.n88 VGND.n75 0.120292
R781 VGND.n88 VGND.n87 0.120292
R782 VGND.n87 VGND.n78 0.120292
R783 VGND.n83 VGND.n78 0.120292
R784 VGND.n83 VGND.n82 0.120292
R785 VGND.n82 VGND.n81 0.120292
R786 VGND.n422 VGND.n421 0.120292
R787 VGND.n423 VGND.n422 0.120292
R788 VGND.n423 VGND.n22 0.120292
R789 VGND.n427 VGND.n22 0.120292
R790 VGND.n428 VGND.n427 0.120292
R791 VGND.n429 VGND.n428 0.120292
R792 VGND.n429 VGND.n19 0.120292
R793 VGND.n433 VGND.n19 0.120292
R794 VGND.n434 VGND.n433 0.120292
R795 VGND.n435 VGND.n434 0.120292
R796 VGND.n435 VGND.n17 0.120292
R797 VGND.n441 VGND.n17 0.120292
R798 VGND.n442 VGND.n441 0.120292
R799 VGND.n443 VGND.n442 0.120292
R800 VGND.n443 VGND.n15 0.120292
R801 VGND.n384 VGND.n333 0.115155
R802 VGND.n404 VGND.n403 0.110794
R803 VGND.n357 VGND.n356 0.110004
R804 VGND.n381 VGND.n337 0.109215
R805 VGND.n356 VGND.n355 0.108082
R806 VGND.n355 VGND.n354 0.105175
R807 VGND.n279 VGND.n246 0.105059
R808 VGND.n359 VGND.n357 0.104833
R809 VGND.n372 VGND.n346 0.104045
R810 VGND.n354 VGND.n353 0.1015
R811 VGND.n353 VGND.n352 0.0997064
R812 VGND.n107 VGND 0.0981562
R813 VGND.n421 VGND 0.0981562
R814 VGND.n352 VGND.n351 0.097941
R815 VGND.n351 VGND.n350 0.0952266
R816 VGND.n337 VGND.n334 0.0946901
R817 VGND.n350 VGND.n349 0.0925543
R818 VGND.n460 VGND.n6 0.0910095
R819 VGND.n349 VGND.n348 0.0892405
R820 VGND.n348 VGND.n347 0.0876212
R821 VGND.n7 VGND.n6 0.0867209
R822 VGND.n457 VGND.n5 0.0867069
R823 VGND.n347 VGND.n346 0.0860263
R824 VGND.n373 VGND.n372 0.0819653
R825 VGND.n345 VGND.n344 0.0807239
R826 VGND.n383 VGND.n382 0.0803467
R827 VGND.n459 VGND.n5 0.0798478
R828 VGND.n458 VGND.n7 0.0787609
R829 VGND.n457 VGND.n456 0.0782778
R830 VGND.n358 VGND.n8 0.0776277
R831 VGND.n344 VGND.n343 0.0771423
R832 VGND.n343 VGND.n342 0.0762299
R833 VGND.n41 VGND 0.0758148
R834 VGND.n342 VGND.n341 0.0738696
R835 VGND.n358 VGND.n6 0.0721983
R836 VGND.n316 VGND.n315 0.0721201
R837 VGND.n461 VGND.n460 0.0720511
R838 VGND.n341 VGND.n340 0.0715432
R839 VGND.n340 VGND.n339 0.0701429
R840 VGND.n382 VGND.n381 0.0683371
R841 VGND.n339 VGND.n338 0.0678759
R842 VGND.n279 VGND.n278 0.0678759
R843 VGND.n333 VGND.n332 0.0675348
R844 VGND.n338 VGND.n337 0.0656408
R845 VGND.n278 VGND.n277 0.0656408
R846 VGND.n277 VGND.n248 0.0638803
R847 VGND.n249 VGND.n248 0.0621319
R848 VGND VGND.n68 0.0603958
R849 VGND.n112 VGND 0.0603958
R850 VGND VGND.n111 0.0603958
R851 VGND VGND.n110 0.0603958
R852 VGND.n81 VGND 0.0603958
R853 VGND.n415 VGND 0.0603958
R854 VGND.n416 VGND 0.0603958
R855 VGND.n417 VGND 0.0603958
R856 VGND.n250 VGND.n249 0.0591207
R857 VGND.n359 VGND.n358 0.0590106
R858 VGND.n251 VGND.n250 0.0582586
R859 VGND.n184 VGND 0.05675
R860 VGND.n244 VGND 0.05675
R861 VGND.n406 VGND 0.05675
R862 VGND.n3 VGND 0.05675
R863 VGND.n4 VGND 0.05675
R864 VGND.n2 VGND 0.05675
R865 VGND.n455 VGND 0.05675
R866 VGND.n336 VGND 0.05675
R867 VGND.n289 VGND 0.05675
R868 VGND.n294 VGND 0.05675
R869 VGND.n282 VGND 0.05675
R870 VGND.n383 VGND.n334 0.0567284
R871 VGND.n332 VGND.n331 0.0561507
R872 VGND.n252 VGND.n251 0.0561507
R873 VGND.n331 VGND.n330 0.0549218
R874 VGND.n253 VGND.n252 0.0549218
R875 VGND.n227 VGND.n226 0.0533169
R876 VGND.n330 VGND.n329 0.0520203
R877 VGND.n254 VGND.n253 0.0520203
R878 VGND.n329 VGND.n328 0.0511757
R879 VGND.n255 VGND.n254 0.0511757
R880 VGND.n228 VGND.n227 0.0509967
R881 VGND.n226 VGND.n155 0.0486419
R882 VGND.n328 VGND.n327 0.0483188
R883 VGND.n256 VGND.n255 0.0483188
R884 VGND.n156 VGND.n155 0.0477973
R885 VGND.n327 VGND.n326 0.0471667
R886 VGND.n257 VGND.n256 0.0471667
R887 VGND.n157 VGND.n156 0.045802
R888 VGND.n326 VGND.n325 0.045202
R889 VGND.n258 VGND.n257 0.045202
R890 VGND.n158 VGND.n157 0.0438333
R891 VGND.n325 VGND.n324 0.0435464
R892 VGND.n259 VGND.n258 0.0435464
R893 VGND.n324 VGND.n323 0.0418907
R894 VGND.n260 VGND.n259 0.0418907
R895 VGND.n159 VGND.n158 0.0418907
R896 VGND.n160 VGND.n159 0.0410629
R897 VGND.n458 VGND.n457 0.0407778
R898 VGND.n402 VGND.n317 0.0407077
R899 VGND.n323 VGND.n322 0.0405327
R900 VGND.n261 VGND.n260 0.0405327
R901 VGND.n161 VGND.n160 0.0385795
R902 VGND.n322 VGND.n321 0.0380817
R903 VGND.n261 VGND.n137 0.0380817
R904 VGND.n321 VGND.n320 0.0364477
R905 VGND.n297 VGND.n137 0.0364477
R906 VGND.n162 VGND.n161 0.0364477
R907 VGND.n163 VGND.n162 0.0356307
R908 VGND.n320 VGND.n319 0.0354026
R909 VGND.n298 VGND.n297 0.0354026
R910 VGND.n112 VGND 0.0343542
R911 VGND.n111 VGND 0.0343542
R912 VGND VGND.n415 0.0343542
R913 VGND VGND.n416 0.0343542
R914 VGND.n281 VGND.n280 0.0341879
R915 VGND.n164 VGND.n163 0.0331797
R916 VGND.n319 VGND.n318 0.0327581
R917 VGND.n299 VGND.n298 0.0327581
R918 VGND.n165 VGND.n164 0.0321558
R919 VGND.n401 VGND.n318 0.0319516
R920 VGND.n300 VGND.n299 0.0319516
R921 VGND.n334 VGND.n333 0.0307768
R922 VGND.n402 VGND.n401 0.0303387
R923 VGND.n301 VGND.n300 0.0303387
R924 VGND.n166 VGND.n165 0.0303387
R925 VGND.n456 VGND.n8 0.0297553
R926 VGND.n229 VGND.n228 0.0292963
R927 VGND.n466 VGND.n0 0.0288333
R928 VGND.n467 VGND.n466 0.0288333
R929 VGND.n167 VGND.n166 0.0279194
R930 VGND.n302 VGND.n301 0.0277436
R931 VGND.n168 VGND.n167 0.0271129
R932 VGND.n303 VGND.n302 0.0269423
R933 VGND.n169 VGND.n168 0.0253397
R934 VGND.n304 VGND.n303 0.0251815
R935 VGND.n170 VGND.n169 0.0237372
R936 VGND.n305 VGND.n304 0.0235892
R937 VGND.n110 VGND 0.0226354
R938 VGND.n417 VGND 0.0226354
R939 VGND.n306 VGND.n305 0.0219968
R940 VGND.n171 VGND.n170 0.0219968
R941 VGND.n307 VGND.n306 0.0204045
R942 VGND.n308 VGND.n307 0.0186962
R943 VGND.n296 VGND.n295 0.0175455
R944 VGND.n309 VGND.n308 0.0171139
R945 VGND.n310 VGND.n309 0.0154371
R946 VGND.n403 VGND.n117 0.0141218
R947 VGND.n311 VGND.n310 0.0139494
R948 VGND.n459 VGND.n458 0.0135435
R949 VGND.n312 VGND.n311 0.0122925
R950 VGND.n313 VGND.n312 0.00993396
R951 VGND.n208 VGND.n171 0.00918938
R952 VGND.n314 VGND.n313 0.0091478
R953 VGND.n315 VGND.n314 0.00757547
R954 VGND.n287 VGND.n119 0.00689301
R955 VGND.n465 VGND.n464 0.0011075
R956 VDPWR.n1 VDPWR.t7 738.801
R957 VDPWR.n1 VDPWR.t6 707.519
R958 VDPWR.n84 VDPWR.t67 667.734
R959 VDPWR.n52 VDPWR.t37 667.734
R960 VDPWR.n124 VDPWR.t51 667.734
R961 VDPWR.n99 VDPWR.t63 666.677
R962 VDPWR.n38 VDPWR.t17 666.677
R963 VDPWR.n4 VDPWR.t47 666.677
R964 VDPWR.t44 VDPWR.t50 624.456
R965 VDPWR.t36 VDPWR.t18 624.456
R966 VDPWR.t66 VDPWR.t48 624.456
R967 VDPWR.n102 VDPWR.n101 604.394
R968 VDPWR.n33 VDPWR.n32 604.394
R969 VDPWR.n142 VDPWR.n141 604.394
R970 VDPWR.t46 VDPWR.t20 556.386
R971 VDPWR.t52 VDPWR.t54 556.386
R972 VDPWR.t40 VDPWR.t16 556.386
R973 VDPWR.t32 VDPWR.t34 556.386
R974 VDPWR.t59 VDPWR.t62 556.386
R975 VDPWR.t70 VDPWR.t68 556.386
R976 VDPWR.n17 VDPWR.t72 414.33
R977 VDPWR.t42 VDPWR.n108 414.33
R978 VDPWR.t0 VDPWR.t4 390.654
R979 VDPWR.t8 VDPWR.t28 390.654
R980 VDPWR.t56 VDPWR.t30 390.654
R981 VDPWR.t50 VDPWR.t3 337.384
R982 VDPWR.t24 VDPWR.t36 337.384
R983 VDPWR.t26 VDPWR.t66 337.384
R984 VDPWR.n82 VDPWR.n72 333.348
R985 VDPWR.n54 VDPWR.n24 333.348
R986 VDPWR.n122 VDPWR.n12 333.348
R987 VDPWR.n68 VDPWR.n67 320.976
R988 VDPWR.n45 VDPWR.n28 320.976
R989 VDPWR.n9 VDPWR.n8 320.976
R990 VDPWR.t4 VDPWR.t23 304.829
R991 VDPWR.t38 VDPWR.t8 304.829
R992 VDPWR.t61 VDPWR.t56 304.829
R993 VDPWR.t72 VDPWR.t52 287.072
R994 VDPWR.t34 VDPWR.t42 287.072
R995 VDPWR.t68 VDPWR.t64 287.072
R996 VDPWR.t23 VDPWR.t2 281.154
R997 VDPWR.t22 VDPWR.t0 281.154
R998 VDPWR.t25 VDPWR.t38 281.154
R999 VDPWR.t28 VDPWR.t39 281.154
R1000 VDPWR.t27 VDPWR.t61 281.154
R1001 VDPWR.t30 VDPWR.t58 281.154
R1002 VDPWR.n109 VDPWR.n17 272.274
R1003 VDPWR.n109 VDPWR 272.274
R1004 VDPWR.n108 VDPWR.n107 272.274
R1005 VDPWR.n107 VDPWR 272.274
R1006 VDPWR.t2 VDPWR.t46 251.559
R1007 VDPWR.t16 VDPWR.t25 251.559
R1008 VDPWR.t62 VDPWR.t27 251.559
R1009 VDPWR.t20 VDPWR.t14 248.599
R1010 VDPWR.t3 VDPWR.t22 248.599
R1011 VDPWR.t54 VDPWR.t44 248.599
R1012 VDPWR.t12 VDPWR.t40 248.599
R1013 VDPWR.t39 VDPWR.t24 248.599
R1014 VDPWR.t18 VDPWR.t32 248.599
R1015 VDPWR.t10 VDPWR.t59 248.599
R1016 VDPWR.t58 VDPWR.t26 248.599
R1017 VDPWR.t48 VDPWR.t70 248.599
R1018 VDPWR.n76 VDPWR.n75 240.522
R1019 VDPWR.n60 VDPWR.n21 240.522
R1020 VDPWR.n116 VDPWR.n115 240.522
R1021 VDPWR.n107 VDPWR.n106 213.119
R1022 VDPWR.n108 VDPWR.n18 213.119
R1023 VDPWR.n110 VDPWR.n109 213.119
R1024 VDPWR.n17 VDPWR.n15 213.119
R1025 VDPWR.n67 VDPWR.t57 113.98
R1026 VDPWR.n28 VDPWR.t9 113.98
R1027 VDPWR.n8 VDPWR.t5 113.98
R1028 VDPWR.t14 VDPWR 91.745
R1029 VDPWR VDPWR.t12 91.745
R1030 VDPWR VDPWR.t10 91.745
R1031 VDPWR.n75 VDPWR.t69 61.9872
R1032 VDPWR.n21 VDPWR.t35 61.9872
R1033 VDPWR.n115 VDPWR.t53 61.9872
R1034 VDPWR.n101 VDPWR.t11 41.5552
R1035 VDPWR.n101 VDPWR.t60 41.5552
R1036 VDPWR.n32 VDPWR.t13 41.5552
R1037 VDPWR.n32 VDPWR.t41 41.5552
R1038 VDPWR.n141 VDPWR.t15 41.5552
R1039 VDPWR.n141 VDPWR.t21 41.5552
R1040 VDPWR.n67 VDPWR.t31 35.4605
R1041 VDPWR.n28 VDPWR.t29 35.4605
R1042 VDPWR.n8 VDPWR.t1 35.4605
R1043 VDPWR.n81 VDPWR.n73 34.6358
R1044 VDPWR.n77 VDPWR.n73 34.6358
R1045 VDPWR.n95 VDPWR.n65 34.6358
R1046 VDPWR.n95 VDPWR.n94 34.6358
R1047 VDPWR.n94 VDPWR.n93 34.6358
R1048 VDPWR.n90 VDPWR.n89 34.6358
R1049 VDPWR.n89 VDPWR.n88 34.6358
R1050 VDPWR.n88 VDPWR.n70 34.6358
R1051 VDPWR.n55 VDPWR.n22 34.6358
R1052 VDPWR.n59 VDPWR.n22 34.6358
R1053 VDPWR.n40 VDPWR.n39 34.6358
R1054 VDPWR.n40 VDPWR.n29 34.6358
R1055 VDPWR.n44 VDPWR.n29 34.6358
R1056 VDPWR.n47 VDPWR.n46 34.6358
R1057 VDPWR.n47 VDPWR.n26 34.6358
R1058 VDPWR.n51 VDPWR.n26 34.6358
R1059 VDPWR.n121 VDPWR.n13 34.6358
R1060 VDPWR.n117 VDPWR.n13 34.6358
R1061 VDPWR.n136 VDPWR.n135 34.6358
R1062 VDPWR.n135 VDPWR.n134 34.6358
R1063 VDPWR.n134 VDPWR.n6 34.6358
R1064 VDPWR.n130 VDPWR.n129 34.6358
R1065 VDPWR.n129 VDPWR.n128 34.6358
R1066 VDPWR.n128 VDPWR.n10 34.6358
R1067 VDPWR.n83 VDPWR.n82 32.0005
R1068 VDPWR.n54 VDPWR.n53 32.0005
R1069 VDPWR.n123 VDPWR.n122 32.0005
R1070 VDPWR.n143 VDPWR.n142 30.7593
R1071 VDPWR.n84 VDPWR.n83 30.4946
R1072 VDPWR.n53 VDPWR.n52 30.4946
R1073 VDPWR.n124 VDPWR.n123 30.4946
R1074 VDPWR.n75 VDPWR.t65 30.1692
R1075 VDPWR.n21 VDPWR.t43 30.1692
R1076 VDPWR.n115 VDPWR.t73 30.1692
R1077 VDPWR.n99 VDPWR.n65 27.4829
R1078 VDPWR.n61 VDPWR.n60 27.4829
R1079 VDPWR.n39 VDPWR.n38 27.4829
R1080 VDPWR.n116 VDPWR.n114 27.4829
R1081 VDPWR.n136 VDPWR.n4 27.4829
R1082 VDPWR.n72 VDPWR.t49 26.5955
R1083 VDPWR.n72 VDPWR.t71 26.5955
R1084 VDPWR.n24 VDPWR.t19 26.5955
R1085 VDPWR.n24 VDPWR.t33 26.5955
R1086 VDPWR.n12 VDPWR.t45 26.5955
R1087 VDPWR.n12 VDPWR.t55 26.5955
R1088 VDPWR.n77 VDPWR.n76 25.6005
R1089 VDPWR.n60 VDPWR.n59 25.6005
R1090 VDPWR.n117 VDPWR.n116 25.6005
R1091 VDPWR.n106 VDPWR.n19 23.7181
R1092 VDPWR.n61 VDPWR.n18 23.7181
R1093 VDPWR.n110 VDPWR.n16 23.7181
R1094 VDPWR.n114 VDPWR.n15 23.7181
R1095 VDPWR.n102 VDPWR.n100 22.9652
R1096 VDPWR.n37 VDPWR.n33 22.9652
R1097 VDPWR.n142 VDPWR.n140 22.9652
R1098 VDPWR.n100 VDPWR.n99 21.8358
R1099 VDPWR.n38 VDPWR.n37 21.8358
R1100 VDPWR.n140 VDPWR.n4 21.8358
R1101 VDPWR.n102 VDPWR.n19 21.4593
R1102 VDPWR.n33 VDPWR.n16 21.4593
R1103 VDPWR.n93 VDPWR.n68 18.4476
R1104 VDPWR.n45 VDPWR.n44 18.4476
R1105 VDPWR.n9 VDPWR.n6 18.4476
R1106 VDPWR.n90 VDPWR.n68 16.1887
R1107 VDPWR.n46 VDPWR.n45 16.1887
R1108 VDPWR.n130 VDPWR.n9 16.1887
R1109 VDPWR.n84 VDPWR.n70 15.0593
R1110 VDPWR.n52 VDPWR.n51 15.0593
R1111 VDPWR.n124 VDPWR.n10 15.0593
R1112 VDPWR.n2 VDPWR.n1 13.3223
R1113 VDPWR.n106 VDPWR.n18 12.8005
R1114 VDPWR.n110 VDPWR.n15 12.8005
R1115 VDPWR.n3 VDPWR 9.73982
R1116 VDPWR.n143 VDPWR.n3 9.61724
R1117 VDPWR.n142 VDPWR.n0 9.3005
R1118 VDPWR.n140 VDPWR.n139 9.3005
R1119 VDPWR.n138 VDPWR.n4 9.3005
R1120 VDPWR.n137 VDPWR.n136 9.3005
R1121 VDPWR.n135 VDPWR.n5 9.3005
R1122 VDPWR.n134 VDPWR.n133 9.3005
R1123 VDPWR.n132 VDPWR.n6 9.3005
R1124 VDPWR.n131 VDPWR.n130 9.3005
R1125 VDPWR.n129 VDPWR.n7 9.3005
R1126 VDPWR.n128 VDPWR.n127 9.3005
R1127 VDPWR.n126 VDPWR.n10 9.3005
R1128 VDPWR.n125 VDPWR.n124 9.3005
R1129 VDPWR.n123 VDPWR.n11 9.3005
R1130 VDPWR.n121 VDPWR.n120 9.3005
R1131 VDPWR.n119 VDPWR.n13 9.3005
R1132 VDPWR.n118 VDPWR.n117 9.3005
R1133 VDPWR.n116 VDPWR.n14 9.3005
R1134 VDPWR.n114 VDPWR.n113 9.3005
R1135 VDPWR.n112 VDPWR.n15 9.3005
R1136 VDPWR.n111 VDPWR.n110 9.3005
R1137 VDPWR.n34 VDPWR.n16 9.3005
R1138 VDPWR.n35 VDPWR.n33 9.3005
R1139 VDPWR.n37 VDPWR.n36 9.3005
R1140 VDPWR.n38 VDPWR.n31 9.3005
R1141 VDPWR.n39 VDPWR.n30 9.3005
R1142 VDPWR.n41 VDPWR.n40 9.3005
R1143 VDPWR.n42 VDPWR.n29 9.3005
R1144 VDPWR.n44 VDPWR.n43 9.3005
R1145 VDPWR.n46 VDPWR.n27 9.3005
R1146 VDPWR.n48 VDPWR.n47 9.3005
R1147 VDPWR.n49 VDPWR.n26 9.3005
R1148 VDPWR.n51 VDPWR.n50 9.3005
R1149 VDPWR.n52 VDPWR.n25 9.3005
R1150 VDPWR.n53 VDPWR.n23 9.3005
R1151 VDPWR.n56 VDPWR.n55 9.3005
R1152 VDPWR.n57 VDPWR.n22 9.3005
R1153 VDPWR.n59 VDPWR.n58 9.3005
R1154 VDPWR.n60 VDPWR.n20 9.3005
R1155 VDPWR.n62 VDPWR.n61 9.3005
R1156 VDPWR.n63 VDPWR.n18 9.3005
R1157 VDPWR.n106 VDPWR.n105 9.3005
R1158 VDPWR.n104 VDPWR.n19 9.3005
R1159 VDPWR.n103 VDPWR.n102 9.3005
R1160 VDPWR.n100 VDPWR.n64 9.3005
R1161 VDPWR.n99 VDPWR.n98 9.3005
R1162 VDPWR.n97 VDPWR.n65 9.3005
R1163 VDPWR.n96 VDPWR.n95 9.3005
R1164 VDPWR.n94 VDPWR.n66 9.3005
R1165 VDPWR.n93 VDPWR.n92 9.3005
R1166 VDPWR.n91 VDPWR.n90 9.3005
R1167 VDPWR.n89 VDPWR.n69 9.3005
R1168 VDPWR.n88 VDPWR.n87 9.3005
R1169 VDPWR.n86 VDPWR.n70 9.3005
R1170 VDPWR.n85 VDPWR.n84 9.3005
R1171 VDPWR.n83 VDPWR.n71 9.3005
R1172 VDPWR.n81 VDPWR.n80 9.3005
R1173 VDPWR.n79 VDPWR.n73 9.3005
R1174 VDPWR.n78 VDPWR.n77 9.3005
R1175 VDPWR.n3 VDPWR.n2 8.39487
R1176 VDPWR.n76 VDPWR.n74 7.4049
R1177 VDPWR.n82 VDPWR.n81 2.63579
R1178 VDPWR.n55 VDPWR.n54 2.63579
R1179 VDPWR.n122 VDPWR.n121 2.63579
R1180 VDPWR.n74 VDPWR 0.156264
R1181 VDPWR.n78 VDPWR.n74 0.144904
R1182 VDPWR.n139 VDPWR.n0 0.120292
R1183 VDPWR.n139 VDPWR.n138 0.120292
R1184 VDPWR.n138 VDPWR.n137 0.120292
R1185 VDPWR.n137 VDPWR.n5 0.120292
R1186 VDPWR.n133 VDPWR.n5 0.120292
R1187 VDPWR.n133 VDPWR.n132 0.120292
R1188 VDPWR.n132 VDPWR.n131 0.120292
R1189 VDPWR.n131 VDPWR.n7 0.120292
R1190 VDPWR.n127 VDPWR.n7 0.120292
R1191 VDPWR.n127 VDPWR.n126 0.120292
R1192 VDPWR.n126 VDPWR.n125 0.120292
R1193 VDPWR.n125 VDPWR.n11 0.120292
R1194 VDPWR.n120 VDPWR.n11 0.120292
R1195 VDPWR.n120 VDPWR.n119 0.120292
R1196 VDPWR.n119 VDPWR.n118 0.120292
R1197 VDPWR.n118 VDPWR.n14 0.120292
R1198 VDPWR.n113 VDPWR.n14 0.120292
R1199 VDPWR.n36 VDPWR.n35 0.120292
R1200 VDPWR.n36 VDPWR.n31 0.120292
R1201 VDPWR.n31 VDPWR.n30 0.120292
R1202 VDPWR.n41 VDPWR.n30 0.120292
R1203 VDPWR.n42 VDPWR.n41 0.120292
R1204 VDPWR.n43 VDPWR.n42 0.120292
R1205 VDPWR.n43 VDPWR.n27 0.120292
R1206 VDPWR.n48 VDPWR.n27 0.120292
R1207 VDPWR.n49 VDPWR.n48 0.120292
R1208 VDPWR.n50 VDPWR.n49 0.120292
R1209 VDPWR.n50 VDPWR.n25 0.120292
R1210 VDPWR.n25 VDPWR.n23 0.120292
R1211 VDPWR.n56 VDPWR.n23 0.120292
R1212 VDPWR.n57 VDPWR.n56 0.120292
R1213 VDPWR.n58 VDPWR.n57 0.120292
R1214 VDPWR.n58 VDPWR.n20 0.120292
R1215 VDPWR.n62 VDPWR.n20 0.120292
R1216 VDPWR.n103 VDPWR.n64 0.120292
R1217 VDPWR.n98 VDPWR.n64 0.120292
R1218 VDPWR.n98 VDPWR.n97 0.120292
R1219 VDPWR.n97 VDPWR.n96 0.120292
R1220 VDPWR.n96 VDPWR.n66 0.120292
R1221 VDPWR.n92 VDPWR.n66 0.120292
R1222 VDPWR.n92 VDPWR.n91 0.120292
R1223 VDPWR.n91 VDPWR.n69 0.120292
R1224 VDPWR.n87 VDPWR.n69 0.120292
R1225 VDPWR.n87 VDPWR.n86 0.120292
R1226 VDPWR.n86 VDPWR.n85 0.120292
R1227 VDPWR.n85 VDPWR.n71 0.120292
R1228 VDPWR.n80 VDPWR.n71 0.120292
R1229 VDPWR.n80 VDPWR.n79 0.120292
R1230 VDPWR.n79 VDPWR.n78 0.120292
R1231 VDPWR VDPWR.n0 0.0981562
R1232 VDPWR.n35 VDPWR 0.0981562
R1233 VDPWR VDPWR.n103 0.0981562
R1234 VDPWR.n113 VDPWR 0.0603958
R1235 VDPWR VDPWR.n112 0.0603958
R1236 VDPWR VDPWR.n111 0.0603958
R1237 VDPWR.n34 VDPWR 0.0603958
R1238 VDPWR VDPWR.n62 0.0603958
R1239 VDPWR.n63 VDPWR 0.0603958
R1240 VDPWR.n105 VDPWR 0.0603958
R1241 VDPWR VDPWR.n104 0.0603958
R1242 VDPWR.n2 VDPWR 0.0496071
R1243 VDPWR.n112 VDPWR 0.0382604
R1244 VDPWR.n111 VDPWR 0.0382604
R1245 VDPWR VDPWR.n63 0.0382604
R1246 VDPWR.n105 VDPWR 0.0382604
R1247 VDPWR VDPWR.n34 0.0226354
R1248 VDPWR.n104 VDPWR 0.0226354
R1249 VDPWR VDPWR.n143 0.0224072
R1250 uo_out[1].n2 uo_out[1].t1 313.104
R1251 uo_out[1].n0 uo_out[1].t2 294.557
R1252 uo_out[1].t0 uo_out[1].n2 265.769
R1253 uo_out[1] uo_out[1].t0 262.318
R1254 uo_out[1].n0 uo_out[1].t3 211.01
R1255 uo_out[1].n1 uo_out[1].n0 152
R1256 uo_out[1].n5 uo_out[1] 12.6752
R1257 uo_out[1].n4 uo_out[1].n1 11.6411
R1258 uo_out[1].n4 uo_out[1].n3 9.3005
R1259 uo_out[1].n3 uo_out[1] 7.17626
R1260 uo_out[1].n3 uo_out[1].n2 4.84898
R1261 uo_out[1].n5 uo_out[1].n4 4.5029
R1262 uo_out[1].n1 uo_out[1] 1.37896
R1263 uo_out[1] uo_out[1].n5 0.0730806
R1264 uo_out[3].n0 uo_out[3].t1 313.104
R1265 uo_out[3].t0 uo_out[3].n0 265.769
R1266 uo_out[3] uo_out[3].t0 262.318
R1267 uo_out[3].n2 uo_out[3] 19.5328
R1268 uo_out[3].n2 uo_out[3].n1 13.8005
R1269 uo_out[3].n1 uo_out[3].n0 7.17626
R1270 uo_out[3].n1 uo_out[3] 4.84898
R1271 uo_out[3] uo_out[3].n2 0.0529194
R1272 uo_out[0].n4 uo_out[0].t1 983.422
R1273 uo_out[0] uo_out[0].t0 455.764
R1274 uo_out[0].n0 uo_out[0].t3 294.557
R1275 uo_out[0].n0 uo_out[0].t2 211.01
R1276 uo_out[0].n1 uo_out[0].n0 152
R1277 uo_out[0].n4 uo_out[0].n3 19.6603
R1278 uo_out[0].n2 uo_out[0].n1 17.6405
R1279 uo_out[0] uo_out[0].n4 10.2862
R1280 uo_out[0].n3 uo_out[0].n2 6.83545
R1281 uo_out[0].n1 uo_out[0] 2.01193
R1282 uo_out[0].n3 uo_out[0] 1.31337
R1283 uo_out[0].n2 uo_out[0] 0.0793043
R1284 uo_out[2].n2 uo_out[2].t1 313.104
R1285 uo_out[2].n0 uo_out[2].t2 294.557
R1286 uo_out[2].t0 uo_out[2].n2 265.769
R1287 uo_out[2] uo_out[2].t0 262.318
R1288 uo_out[2].n0 uo_out[2].t3 211.01
R1289 uo_out[2].n1 uo_out[2].n0 152
R1290 uo_out[2].n5 uo_out[2] 16.2155
R1291 uo_out[2].n4 uo_out[2].n1 11.6311
R1292 uo_out[2].n4 uo_out[2].n3 9.3005
R1293 uo_out[2].n3 uo_out[2] 7.17626
R1294 uo_out[2].n3 uo_out[2].n2 4.84898
R1295 uo_out[2].n5 uo_out[2].n4 4.51042
R1296 uo_out[2].n1 uo_out[2] 1.37896
R1297 uo_out[2] uo_out[2].n5 0.0730806
C0 m2_18496_33616# m1_18496_33616# 2.03601f
C1 m2_5328_26928# m1_5328_26928# 2.03601f
C2 m2_22770_15390# m1_22770_15390# 2.03601f
C3 m2_4416_23566# m1_4416_23566# 2.03601f
C4 m3_11508_25704# m2_11508_25704# 71.142296f
C5 m2_17976_13788# m1_17976_13788# 2.03601f
C6 m2_20662_15338# m1_20662_15338# 2.03601f
C7 m1_24714_26720# m2_24714_26720# 2.03601f
C8 m1_20662_13418# m2_20662_13418# 2.03601f
C9 m1_4708_16904# m2_4708_16904# 2.03601f
C10 m2_10182_17306# m1_10182_17306# 75.185295f
C11 VAPWR VDPWR 19.2978f
C12 m2_17976_11868# m1_17976_11868# 2.03601f
C13 m1_3616_22186# m2_3616_22186# 2.03601f
C14 m1_14954_13098# m2_14954_13098# 2.03601f
C15 m2_9500_32942# m1_9500_32942# 2.03601f
C16 m2_25498_21416# m1_25498_21416# 2.03601f
C17 m1_7588_42050# m2_7588_42050# 2.03601f
C18 m2_11508_25704# m1_11508_25704# 0.11049p
C19 m1_15474_32386# m2_15474_32386# 2.03601f
C20 m2_4416_25486# m1_4416_25486# 2.03601f
C21 m1_7076_29088# m2_7076_29088# 2.03601f
C22 m2_7076_31008# m1_7076_31008# 2.03601f
C23 m1_5328_28848# m2_5328_28848# 2.03601f
C24 m2_6556_14476# m1_6556_14476# 2.03601f
C25 m3_10182_17306# m2_10182_17306# 48.4105f
C26 m2_8978_14462# m1_8978_14462# 2.03601f
C27 m2_21182_32066# m1_21182_32066# 2.03601f
C28 m1_24714_24800# m2_24714_24800# 2.03601f
C29 m2_15474_34306# m1_15474_34306# 2.03601f
C30 m1_24658_19894# m2_24658_19894# 2.03601f
C31 m2_8978_12542# m1_8978_12542# 2.03601f
C32 m1_12384_32154# m2_12384_32154# 2.03601f
C33 m4_11508_25704# m3_11508_25704# 69.3594f
C34 m1_23290_27874# m2_23290_27874# 2.03601f
C35 m1_18496_31696# m2_18496_31696# 2.03601f
C36 m2_4708_18824# m1_4708_18824# 2.03601f
C37 m2_3616_20266# m1_3616_20266# 2.03601f
C38 m2_24658_17974# m1_24658_17974# 2.03601f
C39 m2_11864_13330# m1_11864_13330# 2.03601f
C40 m1_22770_17310# m2_22770_17310# 2.03601f
C41 m2_12384_34074# m1_12384_34074# 2.03601f
C42 m2_9328_42110# m1_9328_42110# 2.03601f
C43 m1_23290_29794# m2_23290_29794# 2.03601f
C44 uo_out[0] VDPWR 2.35179f
C45 m2_25498_23336# m1_25498_23336# 2.03601f
C46 m1_6556_16396# m2_6556_16396# 2.03601f
C47 m2_9500_31022# m1_9500_31022# 2.03601f
C48 m4_10182_17306# m3_10182_17306# 47.1973f
C49 m1_21182_30146# m2_21182_30146# 2.03601f
C50 m2_14954_11178# m1_14954_11178# 2.03601f
C51 m2_11864_11410# m1_11864_11410# 2.03601f
C52 uo_out[0] VGND 4.712002f
C53 uo_out[3] VGND 1.78221f
C54 VAPWR VGND 0.136019p
C55 VDPWR VGND 52.08213f
C56 m4_10182_17306# VGND 9.38538f $ **FLOATING
C57 m4_11508_25704# VGND 7.22411f $ **FLOATING
C58 m3_10182_17306# VGND 10.656599f $ **FLOATING
C59 m3_11508_25704# VGND 8.43615f $ **FLOATING
C60 m2_10182_17306# VGND 9.82879f $ **FLOATING
C61 m2_11508_25704# VGND 7.81967f $ **FLOATING
C62 m1_10182_17306# VGND 25.3587f $ **FLOATING
C63 m1_11508_25704# VGND 30.364098f $ **FLOATING
C64 ring_0/skullfet_inverter_16.A VGND 4.7412f
C65 ring_0/skullfet_inverter_17.A VGND 4.82913f
C66 ring_0/skullfet_inverter_15.A VGND 4.9312f
C67 ring_0/skullfet_inverter_18.A VGND 4.98339f
C68 ring_0/skullfet_inverter_14.A VGND 5.03686f
C69 ring_0/skullfet_inverter_19.A VGND 4.79856f
C70 ring_0/skullfet_inverter_13.A VGND 4.80717f
C71 ring_0/skullfet_inverter_20.A VGND 4.93069f
C72 ring_0/skullfet_inverter_12.A VGND 6.09378f
C73 ring_0/skullfet_inverter_20.Y VGND 5.87809f
C74 ring_0/skullfet_inverter_11.A VGND 5.42552f
C75 ring_0/skullfet_inverter_1.A VGND 5.68046f
C76 ring_0/skullfet_inverter_10.A VGND 5.3549f
C77 ring_0/skullfet_inverter_2.A VGND 5.93376f
C78 ring_0/skullfet_inverter_9.A VGND 4.59492f
C79 ring_0/skullfet_inverter_3.A VGND 5.00062f
C80 ring_0/skullfet_inverter_4.A VGND 5.01468f
C81 ring_0/skullfet_inverter_7.A VGND 4.92037f
C82 ring_0/skullfet_inverter_6.A VGND 4.74003f
C83 ring_0/skullfet_inverter_5.A VGND 4.83065f
C84 skullfet_level_shifter.A VGND 12.6722f
C85 VDPWR.n3 VGND 7.64663f
C86 VAPWR.n66 VGND 2.66987f
C87 VAPWR.n67 VGND 15.3513f
.ends

