* NGSPICE file created from tt_um_oscillating_bones.ext - technology: ihp-sg13g2

.subckt tt_um_oscillating_bones ena clk rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] VGND VDPWR
X0 uo_out[1].t0 a_22205_61585# VGND.t31 VGND.t30 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X1 VDPWR.t40 a_16367_61578# freq_divider_0.sg13g2_dfrbp_2_0.D VDPWR.t0 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X2 VGND.t38 a_17996_61559# a_17075_61640# VGND.t105 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X3 VGND.t50 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_21132_61704# VGND.t49 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X4 a_16707_61717# a_16367_61578# VDPWR.t40 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X5 a_17910_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t28 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X6 a_20876_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t27 VDPWR.t0 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X7 ring_0/inverter_ring_0/skullfet_inverter_19.A ring_0/inverter_ring_0/skullfet_inverter_0.Y VDPWR.t65 VDPWR.t64 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X8 VGND.t82 a_22511_61578# a_22205_61585# VGND.t86 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X9 VGND.t48 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_18252_61704# VGND.t47 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X10 ring_0/inverter_ring_0/skullfet_inverter_6.A ring_0/inverter_ring_0/skullfet_inverter_7.A VDPWR.t15 VDPWR.t14 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X11 VGND.t112 ring_0/inverter_ring_0/skullfet_inverter_13.A ring_0/inverter_ring_0/skullfet_inverter_12.A VGND.t111 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X12 VDPWR.t23 a_20876_61559# a_19955_61640# VDPWR.t0 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X13 a_23109_61717# a_22851_61717# VGND.t35 VGND.t34 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X14 a_24054_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t16 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X15 VGND.t72 ring_0/inverter_ring_0/skullfet_inverter_17.A ring_0/inverter_ring_0/skullfet_inverter_16.A VGND.t71 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X16 VGND.t46 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_16801_61717# VGND.t45 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X17 a_20876_61559# a_19947_61366# a_20747_61559# VGND.t76 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X18 ring_0/inverter_ring_0/skullfet_inverter_12.A ring_0/inverter_ring_0/skullfet_inverter_13.A VDPWR.t73 VDPWR.t72 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X19 VDPWR.t54 a_22511_61578# freq_divider_0.sg13g2_dfrbp_2_2.D VDPWR.t0 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X20 a_23211_61366# a_23350_61250# a_23663_61281# VDPWR.t0 sg13_lv_pmos ad=0.3864p pd=2.93u as=0.43102p ps=2.145u w=1.12u l=0.13u
X21 a_23211_61366# a_23350_61250# a_23668_61632# VGND.t8 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.43315p ps=2.205u w=0.74u l=0.13u
X22 VGND.t80 ring_0/inverter_ring_0/skullfet_inverter_9.A ring_0/inverter_ring_0/skullfet_inverter_8.A VGND.t79 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X23 ring_0/inverter_ring_0/skullfet_inverter_11.A ring_0/inverter_ring_0/skullfet_inverter_12.A VDPWR.t43 VDPWR.t42 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X24 VDPWR.t66 freq_divider_0.sg13g2_dfrbp_2_2.D a_24054_61326# VDPWR.t0 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X25 a_22851_61717# a_22511_61578# VDPWR.t54 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X26 a_23161_61402# a_22851_61717# a_23039_61402# VDPWR.t0 sg13_lv_pmos ad=52.5f pd=0.67u as=0.25605p ps=1.935u w=0.42u l=0.13u
X27 VDPWR.t38 a_16367_61578# a_16061_61585# VDPWR.t0 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X28 a_17996_61559# a_17067_61366# a_17867_61559# VGND.t107 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X29 freq_divider_0.sg13g2_dfrbp_2_1.D a_19247_61578# VDPWR.t74 VDPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X30 VDPWR.t3 a_21777_61520# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t0 sg13_lv_pmos ad=0.4657p pd=2.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X31 a_22945_61717# a_22511_61578# a_22851_61717# VGND.t85 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X32 VGND.t44 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_24396_61704# VGND.t43 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X33 VDPWR.t52 a_22511_61578# a_22205_61585# VDPWR.t0 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X34 ring_0/inverter_ring_0/skullfet_inverter_3.A ring_0/inverter_ring_0/skullfet_inverter_4.A VDPWR.t63 VDPWR.t62 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X35 a_24396_61704# a_23219_61640# a_24011_61559# VGND.t21 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X36 a_21856_61617# a_21980_61316# VDPWR.t3 VDPWR.t0 sg13_lv_pmos ad=0.2442p pd=2.06u as=0.4657p ps=2.54u w=0.66u l=0.13u
X37 uo_out[2].t0 a_18941_61585# VGND.t3 VGND.t2 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X38 ring_0/inverter_ring_0/skullfet_inverter_17.A ring_0/inverter_ring_0/skullfet_inverter_18.A VDPWR.t47 VDPWR.t46 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X39 VGND.t33 ring_0/inverter_ring_0/skullfet_inverter_14.A ring_0/inverter_ring_0/skullfet_inverter_13.A VGND.t32 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X40 uo_out[2].t1 a_18941_61585# VDPWR.t2 VDPWR.t0 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X41 VGND.t57 ring_0/inverter_ring_0/skullfet_inverter_2.A ring_0/inverter_ring_0/skullfet_inverter_1.A VGND.t56 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X42 a_19247_61578# a_19947_61366# a_19897_61402# VDPWR.t0 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X43 ring_0/inverter_ring_0/skullfet_inverter_4.A ring_0/inverter_ring_0/skullfet_inverter_5.A VDPWR.t9 VDPWR.t8 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X44 VGND.t90 ring_0/inverter_ring_0/skullfet_inverter_11.A ring_0/inverter_ring_0/skullfet_inverter_10.A VGND.t89 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X45 VDPWR.t1 a_18941_61585# uo_out[2].t1 VDPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X46 VGND.t102 ring_0/inverter_ring_0/skullfet_inverter_0.A ring_0/inverter_ring_0/skullfet_inverter_0.Y VGND.t101 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X47 a_20876_61559# a_19947_61366# a_20790_61326# VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X48 a_18106_61326# a_17206_61250# a_17996_61559# VDPWR.t0 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X49 VGND.t5 ring_0/inverter_ring_0/skullfet_inverter_3.A ring_0/inverter_ring_0/skullfet_inverter_2.A VGND.t4 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X50 VGND.t27 ring_0/inverter_ring_0/skullfet_inverter_16.A uo_out[0].t0 VGND.t26 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X51 ring_0/inverter_ring_0/skullfet_inverter_18.A ring_0/inverter_ring_0/skullfet_inverter_19.A VDPWR.t57 VDPWR.t56 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X52 a_19947_61366# a_20086_61250# a_20399_61281# VDPWR.t0 sg13_lv_pmos ad=0.3864p pd=2.93u as=0.43102p ps=2.145u w=1.12u l=0.13u
X53 ring_0/inverter_ring_0/skullfet_inverter_9.A ring_0/inverter_ring_0/skullfet_inverter_10.A VDPWR.t37 VDPWR.t36 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X54 VGND.t84 a_22511_61578# freq_divider_0.sg13g2_dfrbp_2_2.D VGND.t83 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X55 VGND.t12 uo_out[0].t2 ring_0/inverter_ring_0/skullfet_inverter_14.A VGND.t11 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X56 VGND.t29 a_22205_61585# uo_out[1].t0 VGND.t28 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X57 a_19681_61717# a_19247_61578# a_19587_61717# VGND.t118 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X58 a_17996_61559# a_17067_61366# a_17910_61326# VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X59 a_19955_61640# a_20086_61250# a_19247_61578# VDPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X60 a_20986_61326# a_20086_61250# a_20876_61559# VDPWR.t0 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X61 a_16895_61402# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_16707_61717# VDPWR.t0 sg13_lv_pmos ad=0.25605p pd=1.935u as=79.8f ps=0.8u w=0.42u l=0.13u
X62 a_24140_61559# a_23211_61366# a_24054_61326# VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X63 a_17067_61366# a_17206_61250# a_17519_61281# VDPWR.t0 sg13_lv_pmos ad=0.3864p pd=2.93u as=0.43102p ps=2.145u w=1.12u l=0.13u
X64 a_23039_61402# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_22851_61717# VDPWR.t0 sg13_lv_pmos ad=0.25605p pd=1.935u as=79.8f ps=0.8u w=0.42u l=0.13u
X65 a_17067_61366# a_17206_61250# a_17524_61632# VGND.t99 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.43315p ps=2.205u w=0.74u l=0.13u
X66 VDPWR.t35 freq_divider_0.sg13g2_dfrbp_2_0.D a_17910_61326# VDPWR.t0 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X67 freq_divider_0.sg13g2_dfrbp_2_1.D a_19247_61578# VGND.t114 VGND.t117 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X68 a_21132_61704# a_19955_61640# a_20747_61559# VGND.t108 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X69 a_17910_61326# a_17206_61250# a_17996_61559# VGND.t110 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X70 a_19845_61717# a_20086_61250# a_19247_61578# VGND.t17 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X71 a_16965_61717# a_16707_61717# VGND.t46 VGND.t45 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X72 a_19897_61402# a_19587_61717# a_19775_61402# VDPWR.t0 sg13_lv_pmos ad=52.5f pd=0.67u as=0.25605p ps=1.935u w=0.42u l=0.13u
X73 a_20790_61326# a_20086_61250# a_20876_61559# VGND.t16 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X74 a_18252_61704# a_17075_61640# a_17867_61559# VGND.t54 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X75 VGND.t116 a_19247_61578# freq_divider_0.sg13g2_dfrbp_2_1.D VGND.t115 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X76 VGND.t1 a_18941_61585# uo_out[2].t0 VGND.t0 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X77 a_24140_61559# a_23211_61366# a_24011_61559# VGND.t68 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X78 a_16965_61717# a_17206_61250# a_16367_61578# VGND.t109 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X79 VGND.t114 a_19247_61578# a_18941_61585# VGND.t113 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X80 a_17996_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t25 VDPWR.t0 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X81 VDPWR.t27 a_19955_61640# a_20986_61326# VDPWR.t0 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X82 a_20790_61326# freq_divider_0.sg13g2_dfrbp_2_1.D a_21529_61717# VGND.t53 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X83 VDPWR.t28 a_17996_61559# a_17075_61640# VDPWR.t0 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X84 VGND.t98 ring_0/inverter_ring_0/skullfet_inverter_0.Y ring_0/inverter_ring_0/skullfet_inverter_19.A VGND.t97 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X85 a_24140_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t13 VDPWR.t0 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X86 ring_0/inverter_ring_0/skullfet_inverter_5.A ring_0/inverter_ring_0/skullfet_inverter_6.A VDPWR.t11 VDPWR.t10 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X87 VDPWR.t75 a_19247_61578# freq_divider_0.sg13g2_dfrbp_2_1.D VDPWR.t0 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X88 VGND.t78 ring_0/inverter_ring_0/skullfet_inverter_8.A ring_0/inverter_ring_0/skullfet_inverter_7.A VGND.t77 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X89 a_20399_61281# uo_out[1].t2 a_20086_61250# VDPWR.t0 sg13_lv_pmos ad=0.43102p pd=2.145u as=0.3808p ps=2.92u w=1.12u l=0.13u
X90 VDPWR.t16 a_24140_61559# a_23219_61640# VDPWR.t0 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X91 a_23219_61640# a_23350_61250# a_22511_61578# VDPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X92 VDPWR.t25 a_17075_61640# a_18106_61326# VDPWR.t0 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X93 a_19587_61717# a_19247_61578# VDPWR.t75 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X94 VGND.t52 ring_0/inverter_ring_0/skullfet_inverter_1.A ring_0/inverter_ring_0/skullfet_inverter_0.A VGND.t51 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X95 ring_0/inverter_ring_0/skullfet_inverter_10.A ring_0/inverter_ring_0/skullfet_inverter_11.A VDPWR.t59 VDPWR.t58 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X96 VDPWR.t20 a_22205_61585# uo_out[1].t1 VDPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X97 a_17519_61281# uo_out[2].t2 a_17206_61250# VDPWR.t0 sg13_lv_pmos ad=0.43102p pd=2.145u as=0.3808p ps=2.92u w=1.12u l=0.13u
X98 VGND.t70 ring_0/inverter_ring_0/skullfet_inverter_12.A ring_0/inverter_ring_0/skullfet_inverter_11.A VGND.t69 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X99 a_23109_61717# a_23350_61250# a_22511_61578# VGND.t7 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X100 ring_0/inverter_ring_0/skullfet_inverter_0.A ring_0/inverter_ring_0/skullfet_inverter_1.A VDPWR.t30 VDPWR.t29 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X101 ring_0/inverter_ring_0/skullfet_inverter_16.A ring_0/inverter_ring_0/skullfet_inverter_17.A VDPWR.t45 VDPWR.t44 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X102 a_21980_61316# a_21980_61316# VGND.t10 VGND.t20 sg13_lv_nmos ad=0.111p pd=1.34u as=0.20432p ps=1.585u w=0.3u l=0.13u
X103 VGND.t42 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_19681_61717# VGND.t41 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X104 ring_0/inverter_ring_0/skullfet_inverter_2.A ring_0/inverter_ring_0/skullfet_inverter_3.A VDPWR.t5 VDPWR.t4 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X105 uo_out[0].t1 ring_0/inverter_ring_0/skullfet_inverter_16.A VDPWR.t18 VDPWR.t17 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X106 a_21529_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t40 VGND.t39 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X107 VGND.t40 a_20876_61559# a_19955_61640# VGND.t103 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X108 uo_out[3].t0 a_16061_61585# VGND.t94 VGND.t93 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X109 a_20404_61632# uo_out[1].t2 a_20086_61250# VGND.t15 sg13_lv_nmos ad=0.43315p pd=2.205u as=0.2516p ps=2.16u w=0.74u l=0.13u
X110 VGND.t10 a_21856_61617# a_21777_61520# VGND.t9 sg13_lv_nmos ad=0.20432p pd=1.585u as=0.27427p ps=2.28u w=0.795u l=0.13u
X111 a_16367_61578# a_17067_61366# a_17017_61402# VDPWR.t0 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X112 ring_0/inverter_ring_0/skullfet_inverter_14.A uo_out[0].t2 VDPWR.t7 VDPWR.t6 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X113 VGND.t96 ring_0/inverter_ring_0/skullfet_inverter_4.A ring_0/inverter_ring_0/skullfet_inverter_3.A VGND.t95 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X114 VDPWR.t13 a_23219_61640# a_24250_61326# VDPWR.t0 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X115 a_24250_61326# a_23350_61250# a_24140_61559# VDPWR.t0 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X116 a_20790_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t23 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X117 a_24054_61326# freq_divider_0.sg13g2_dfrbp_2_2.D a_24793_61717# VGND.t100 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X118 a_22511_61578# a_23211_61366# a_23219_61640# VGND.t67 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X119 a_18649_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t38 VGND.t37 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X120 freq_divider_0.sg13g2_dfrbp_2_0.D a_16367_61578# VDPWR.t38 VDPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X121 a_17524_61632# uo_out[2].t2 a_17206_61250# VGND.t99 sg13_lv_nmos ad=0.43315p pd=2.205u as=0.2516p ps=2.16u w=0.74u l=0.13u
X122 VDPWR.t74 a_19247_61578# a_18941_61585# VDPWR.t0 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X123 VGND.t23 ring_0/inverter_ring_0/skullfet_inverter_7.A ring_0/inverter_ring_0/skullfet_inverter_6.A VGND.t22 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X124 a_24793_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t25 VGND.t36 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X125 a_17075_61640# a_17206_61250# a_16367_61578# VDPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X126 uo_out[3].t1 a_16061_61585# VDPWR.t61 VDPWR.t0 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X127 a_24054_61326# a_23350_61250# a_24140_61559# VGND.t6 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X128 VDPWR.t60 a_16061_61585# uo_out[3].t1 VDPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X129 a_22511_61578# a_23211_61366# a_23161_61402# VDPWR.t0 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X130 ring_0/inverter_ring_0/skullfet_inverter_8.A ring_0/inverter_ring_0/skullfet_inverter_9.A VDPWR.t51 VDPWR.t50 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X131 uo_out[1].t1 a_22205_61585# VDPWR.t19 VDPWR.t0 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X132 ring_0/inverter_ring_0/skullfet_inverter_7.A ring_0/inverter_ring_0/skullfet_inverter_8.A VDPWR.t49 VDPWR.t48 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X133 VGND.t60 ring_0/inverter_ring_0/skullfet_inverter_10.A ring_0/inverter_ring_0/skullfet_inverter_9.A VGND.t59 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X134 VGND.t25 a_24140_61559# a_23219_61640# VGND.t24 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X135 a_23668_61632# uo_out[0].t3 a_23350_61250# VGND.t8 sg13_lv_nmos ad=0.43315p pd=2.205u as=0.2516p ps=2.16u w=0.74u l=0.13u
X136 freq_divider_0.sg13g2_dfrbp_2_2.D a_22511_61578# VDPWR.t52 VDPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X137 a_16801_61717# a_16367_61578# a_16707_61717# VGND.t66 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X138 a_19247_61578# a_19947_61366# a_19955_61640# VGND.t75 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X139 ring_0/inverter_ring_0/skullfet_inverter_1.A ring_0/inverter_ring_0/skullfet_inverter_2.A VDPWR.t34 VDPWR.t33 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X140 ring_0/inverter_ring_0/skullfet_inverter_13.A ring_0/inverter_ring_0/skullfet_inverter_14.A VDPWR.t22 VDPWR.t21 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X141 a_19775_61402# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_19587_61717# VDPWR.t0 sg13_lv_pmos ad=0.25605p pd=1.935u as=79.8f ps=0.8u w=0.42u l=0.13u
X142 ring_0/inverter_ring_0/skullfet_inverter_0.Y ring_0/inverter_ring_0/skullfet_inverter_0.A VDPWR.t68 VDPWR.t67 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X143 freq_divider_0.sg13g2_dfrbp_2_0.D a_16367_61578# VGND.t62 VGND.t65 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X144 a_17910_61326# freq_divider_0.sg13g2_dfrbp_2_0.D a_18649_61717# VGND.t58 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X145 a_16367_61578# a_17067_61366# a_17075_61640# VGND.t106 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X146 VGND.t35 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_22945_61717# VGND.t34 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X147 a_17017_61402# a_16707_61717# a_16895_61402# VDPWR.t0 sg13_lv_pmos ad=52.5f pd=0.67u as=0.25605p ps=1.935u w=0.42u l=0.13u
X148 VGND.t74 ring_0/inverter_ring_0/skullfet_inverter_18.A ring_0/inverter_ring_0/skullfet_inverter_17.A VGND.t73 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X149 VGND.t64 a_16367_61578# freq_divider_0.sg13g2_dfrbp_2_0.D VGND.t63 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X150 VGND.t19 ring_0/inverter_ring_0/skullfet_inverter_6.A ring_0/inverter_ring_0/skullfet_inverter_5.A VGND.t18 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X151 VGND.t92 a_16061_61585# uo_out[3].t0 VGND.t91 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X152 a_19845_61717# a_19587_61717# VGND.t42 VGND.t41 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X153 VGND.t14 ring_0/inverter_ring_0/skullfet_inverter_5.A ring_0/inverter_ring_0/skullfet_inverter_4.A VGND.t13 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X154 VGND.t62 a_16367_61578# a_16061_61585# VGND.t61 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X155 a_23663_61281# uo_out[0].t3 a_23350_61250# VDPWR.t0 sg13_lv_pmos ad=0.43102p pd=2.145u as=0.3808p ps=2.92u w=1.12u l=0.13u
X156 a_19947_61366# a_20086_61250# a_20404_61632# VGND.t15 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.43315p ps=2.205u w=0.74u l=0.13u
X157 VGND.t88 ring_0/inverter_ring_0/skullfet_inverter_19.A ring_0/inverter_ring_0/skullfet_inverter_18.A VGND.t87 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X158 VDPWR.t31 freq_divider_0.sg13g2_dfrbp_2_1.D a_20790_61326# VDPWR.t0 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X159 freq_divider_0.sg13g2_dfrbp_2_2.D a_22511_61578# VGND.t82 VGND.t81 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
R0 VGND.n202 VGND.n59 36337.9
R1 VGND.n210 VGND.n111 26006.8
R2 VGND.n349 VGND.n111 20289.4
R3 VGND.t95 VGND.n160 19416.2
R4 VGND.n472 VGND.n471 17662.9
R5 VGND.n194 VGND.n70 15262.5
R6 VGND.n202 VGND.n111 12285.4
R7 VGND.n61 VGND.n59 12285.4
R8 VGND.n471 VGND.n470 12279.6
R9 VGND.n200 VGND.t18 12039.2
R10 VGND.t22 VGND.n63 10402.1
R11 VGND.n285 VGND.n278 10052.7
R12 VGND.n473 VGND.n472 10011.4
R13 VGND.n159 VGND.n158 9840.79
R14 VGND.n201 VGND.n61 9066.9
R15 VGND.n269 VGND.n200 7844.55
R16 VGND.n210 VGND.n204 7498.6
R17 VGND.n199 VGND.n198 7474.99
R18 VGND.n158 VGND.n155 7291.79
R19 VGND.n194 VGND.t13 7169.54
R20 VGND.n476 VGND.n65 6899.39
R21 VGND.n480 VGND.n60 6851.13
R22 VGND.n69 VGND.n65 6429.23
R23 VGND.n269 VGND.t4 6051.63
R24 VGND.n203 VGND.n202 6014.02
R25 VGND.n470 VGND.n469 5872.62
R26 VGND.n204 VGND.n203 5699.78
R27 VGND.n470 VGND.n69 5321.16
R28 VGND.n195 VGND.n194 5298.87
R29 VGND.n482 VGND.n481 4953.11
R30 VGND.n472 VGND.n69 4950.06
R31 VGND.n268 VGND.n267 4945.91
R32 VGND.n295 VGND.n155 3511.45
R33 VGND.n158 VGND.n157 3475.34
R34 VGND.n280 VGND.n275 3284.18
R35 VGND.n470 VGND.n71 3154.9
R36 VGND.n200 VGND.n199 3153.12
R37 VGND.n286 VGND.n285 2376.2
R38 VGND.n269 VGND.n157 2220.92
R39 VGND.n474 VGND.n473 2091.57
R40 VGND.n478 VGND.n63 1946.24
R41 VGND.n203 VGND.n201 1880.71
R42 VGND.n160 VGND.n70 1835.32
R43 VGND.n74 VGND.n71 1763.01
R44 VGND.n269 VGND.n201 1734.38
R45 VGND.n200 VGND.n63 1470.05
R46 VGND.n287 VGND.t101 1368.89
R47 VGND.t87 VGND.n280 1347.06
R48 VGND.n280 VGND.t97 1194.61
R49 VGND.t13 VGND.n193 1123.79
R50 VGND.n471 VGND.n70 1061.65
R51 VGND.n287 VGND.n275 977.779
R52 VGND.n60 VGND.t111 964.287
R53 VGND.n269 VGND.n159 905.553
R54 VGND.t111 VGND.n59 876.317
R55 VGND.n480 VGND.n61 837.723
R56 VGND.n279 VGND.n155 814.62
R57 VGND.n239 VGND.n236 744.615
R58 VGND.n491 VGND.n5 744.615
R59 VGND.n53 VGND.n52 744.615
R60 VGND.n209 VGND.t11 675.663
R61 VGND.n198 VGND.t4 656.004
R62 VGND.n469 VGND.t18 656.004
R63 VGND.n199 VGND.t95 615.229
R64 VGND.n159 VGND.n154 608.424
R65 VGND.n350 VGND.n59 575.212
R66 VGND.n199 VGND.n195 498.868
R67 VGND.n239 VGND.t34 480
R68 VGND.n491 VGND.t41 480
R69 VGND.n52 VGND.t45 480
R70 VGND.n475 VGND.t79 455.887
R71 VGND.n74 VGND.t22 427.755
R72 VGND.n269 VGND.n268 402.269
R73 VGND.n481 VGND.n480 395.865
R74 VGND.n269 VGND.n204 392.892
R75 VGND.t32 VGND.n349 372.399
R76 VGND.n286 VGND.n275 344.149
R77 VGND.t97 VGND.n278 335.173
R78 VGND.n68 VGND.t79 330.428
R79 VGND.n295 VGND.t71 318.406
R80 VGND.n349 VGND.n348 307.757
R81 VGND.n160 VGND.n157 278.079
R82 VGND.n235 VGND.t83 260.005
R83 VGND.n16 VGND.t115 260.005
R84 VGND.t63 VGND.n54 260.005
R85 VGND.t81 VGND.n233 234.738
R86 VGND.t117 VGND.n14 234.738
R87 VGND.n56 VGND.t65 234.738
R88 VGND.n246 VGND.t86 232.869
R89 VGND.n25 VGND.t113 232.869
R90 VGND.t61 VGND.n43 232.869
R91 VGND.t56 VGND.n154 231.615
R92 VGND.t9 VGND.n228 228.233
R93 VGND.n279 VGND.t51 227.947
R94 VGND.n201 VGND.n63 226.054
R95 VGND.n253 VGND.t103 200.339
R96 VGND.n31 VGND.t105 200.339
R97 VGND.n215 VGND.t24 200.339
R98 VGND.n251 VGND.t53 195.942
R99 VGND.n12 VGND.t58 194.969
R100 VGND.n479 VGND.n478 194.851
R101 VGND.n250 VGND.t28 185.124
R102 VGND.n29 VGND.t0 185.124
R103 VGND.t91 VGND.n41 185.124
R104 VGND.t30 VGND.n231 184.825
R105 VGND.t2 VGND.n12 184.825
R106 VGND.n267 VGND.t100 180.052
R107 VGND.n231 VGND.t20 172.145
R108 VGND.n482 VGND.t93 169.907
R109 VGND.n285 VGND.t73 164.255
R110 VGND.t108 VGND.t49 159.763
R111 VGND.t54 VGND.t47 159.763
R112 VGND.t21 VGND.t43 159.763
R113 VGND.t76 VGND.n224 156.929
R114 VGND.t107 VGND.n9 156.929
R115 VGND.t68 VGND.n212 156.929
R116 VGND.n257 VGND.t16 154.614
R117 VGND.n35 VGND.t110 154.614
R118 VGND.n218 VGND.t6 154.614
R119 VGND.n71 VGND.n65 151.276
R120 VGND.t39 VGND.n226 149.62
R121 VGND.t37 VGND.n11 149.62
R122 VGND.t36 VGND.n214 149.62
R123 VGND.t34 VGND.t67 138.463
R124 VGND.t41 VGND.t75 138.463
R125 VGND.t45 VGND.t106 138.463
R126 VGND.n268 VGND.t26 132.323
R127 VGND.n478 VGND.t77 128.216
R128 VGND.n481 VGND.n59 122.921
R129 VGND.t101 VGND.n286 113.026
R130 VGND.n236 VGND.t85 110.237
R131 VGND.t118 VGND.n5 110.237
R132 VGND.t66 VGND.n53 110.237
R133 VGND.n224 VGND.n5 106.212
R134 VGND.n53 VGND.n9 106.212
R135 VGND.n236 VGND.n212 106.212
R136 VGND.t16 VGND.n256 100.478
R137 VGND.t110 VGND.n34 100.478
R138 VGND.t6 VGND.n217 100.478
R139 VGND.n257 VGND.t76 99.7516
R140 VGND.n35 VGND.t107 99.7516
R141 VGND.n218 VGND.t68 99.7516
R142 VGND.n473 VGND.n68 95.8456
R143 VGND.t77 VGND.n477 95.5275
R144 VGND.n253 VGND.t39 93.8297
R145 VGND.n31 VGND.t37 93.8297
R146 VGND.n215 VGND.t36 93.8297
R147 VGND.t20 VGND.n228 86.222
R148 VGND.n295 VGND.n154 84.6642
R149 VGND.n477 VGND.n476 83.8532
R150 VGND.n256 VGND.t108 75.5501
R151 VGND.n34 VGND.t54 75.5501
R152 VGND.n217 VGND.t21 75.5501
R153 VGND.t8 VGND.t7 73.8467
R154 VGND.t15 VGND.t17 73.8467
R155 VGND.t99 VGND.t109 73.8467
R156 VGND.n250 VGND.t30 73.5423
R157 VGND.n29 VGND.t2 73.5423
R158 VGND.t93 VGND.n41 73.5423
R159 VGND.t28 VGND.n246 73.244
R160 VGND.t0 VGND.n25 73.244
R161 VGND.n43 VGND.t91 73.244
R162 VGND.n294 VGND.t51 72.396
R163 VGND.n348 VGND.t11 65.0575
R164 VGND.n350 VGND.t32 63.8663
R165 VGND.n480 VGND.t69 63.5677
R166 VGND.t53 VGND.n226 63.3986
R167 VGND.t58 VGND.n11 63.3986
R168 VGND.n214 VGND.t100 63.3986
R169 VGND.t24 VGND.n213 59.0031
R170 VGND.t103 VGND.n225 59.0031
R171 VGND.t105 VGND.n10 59.0031
R172 VGND.n478 VGND.t89 55.0827
R173 VGND.n270 VGND.t56 51.425
R174 VGND.n206 VGND.t71 51.1311
R175 VGND.t85 VGND.n235 48.4827
R176 VGND.n16 VGND.t118 48.4827
R177 VGND.n54 VGND.t66 48.4827
R178 VGND.t69 VGND.n479 47.9255
R179 VGND.n475 VGND.t59 47.7166
R180 VGND.n475 VGND.n66 44.7738
R181 VGND.n296 VGND.t73 44.7032
R182 VGND.t26 VGND.n210 42.4247
R183 VGND.n66 VGND.t89 41.6077
R184 VGND.n284 VGND.t87 38.7252
R185 VGND.t49 VGND.n225 38.7147
R186 VGND.t47 VGND.n10 38.7147
R187 VGND.t43 VGND.n213 38.7147
R188 VGND.n285 VGND.n279 36.6123
R189 VGND.t59 VGND.n474 36.1063
R190 VGND.n251 VGND.t9 31.1079
R191 VGND.t86 VGND.n233 28.3754
R192 VGND.t113 VGND.n14 28.3754
R193 VGND.n56 VGND.t61 28.3754
R194 VGND.n234 VGND.t81 27.8464
R195 VGND.n15 VGND.t117 27.8464
R196 VGND.t65 VGND.n55 27.8464
R197 VGND.t67 VGND.t8 24.6159
R198 VGND.t75 VGND.t15 24.6159
R199 VGND.t106 VGND.t99 24.6159
R200 VGND.n295 VGND.n294 22.6588
R201 VGND.n210 VGND.n209 22.6333
R202 VGND.n476 VGND.n475 18.8055
R203 VGND.n293 VGND.n292 18.1658
R204 VGND.n272 VGND.n271 18.1658
R205 VGND.n88 VGND.n62 18.1658
R206 VGND.n397 VGND.n396 18.1658
R207 VGND.n77 VGND.n64 18.1658
R208 VGND.n76 VGND.n75 18.1658
R209 VGND.n468 VGND.n467 18.1658
R210 VGND.n193 VGND.n192 18.1658
R211 VGND.n162 VGND.n161 18.1658
R212 VGND.n452 VGND.n451 18.1658
R213 VGND.n87 VGND.n67 18.1658
R214 VGND.n208 VGND.n207 18.1658
R215 VGND.n298 VGND.n297 18.1658
R216 VGND.n283 VGND.n282 18.1658
R217 VGND.n277 VGND.n276 18.1658
R218 VGND.n205 VGND.n141 18.1658
R219 VGND.n347 VGND.n346 18.1658
R220 VGND.n352 VGND.n351 18.1658
R221 VGND.n378 VGND.n377 18.1658
R222 VGND.n197 VGND.n196 18.1658
R223 VGND.n289 VGND.n288 18.1658
R224 VGND.n260 VGND.n257 18.0261
R225 VGND.n489 VGND.n35 18.0261
R226 VGND.n266 VGND.n218 18.0261
R227 VGND.t83 VGND.n234 17.5282
R228 VGND.t115 VGND.n15 17.5282
R229 VGND.n55 VGND.t63 17.5282
R230 VGND.n216 VGND.t25 17.2928
R231 VGND.n36 VGND.t48 17.2395
R232 VGND.n258 VGND.t50 17.2395
R233 VGND.n219 VGND.t44 17.2395
R234 VGND.n47 VGND.t64 17.2297
R235 VGND.n21 VGND.t116 17.2297
R236 VGND.n242 VGND.t84 17.2297
R237 VGND.n40 VGND.t46 17.2268
R238 VGND.n32 VGND.t38 17.2268
R239 VGND.n19 VGND.t42 17.2268
R240 VGND.n254 VGND.t40 17.2268
R241 VGND.n223 VGND.t35 17.2268
R242 VGND.n408 VGND.t62 17.212
R243 VGND.n23 VGND.t114 17.212
R244 VGND.n244 VGND.t82 17.212
R245 VGND.n57 VGND.t94 17.2025
R246 VGND.n27 VGND.t3 17.2025
R247 VGND.n248 VGND.t31 17.2025
R248 VGND.n229 VGND.t10 17.174
R249 VGND.n293 VGND.t52 17.0362
R250 VGND.n271 VGND.t57 17.0362
R251 VGND.n62 VGND.t70 17.0362
R252 VGND.n396 VGND.t90 17.0362
R253 VGND.n64 VGND.t78 17.0362
R254 VGND.n75 VGND.t23 17.0362
R255 VGND.n468 VGND.t19 17.0362
R256 VGND.n193 VGND.t14 17.0362
R257 VGND.n161 VGND.t96 17.0362
R258 VGND.n451 VGND.t80 17.0362
R259 VGND.n67 VGND.t60 17.0362
R260 VGND.n208 VGND.t27 17.0362
R261 VGND.n297 VGND.t74 17.0362
R262 VGND.n283 VGND.t88 17.0362
R263 VGND.n277 VGND.t98 17.0362
R264 VGND.n205 VGND.t72 17.0362
R265 VGND.n347 VGND.t12 17.0362
R266 VGND.n351 VGND.t33 17.0362
R267 VGND.n377 VGND.t112 17.0362
R268 VGND.n197 VGND.t5 17.0362
R269 VGND.n288 VGND.t102 17.0362
R270 VGND.n267 VGND.n266 17.0005
R271 VGND.n266 VGND.n214 17.0005
R272 VGND.n266 VGND.n215 17.0005
R273 VGND.n261 VGND.n260 17.0005
R274 VGND.n260 VGND.n233 17.0005
R275 VGND.n260 VGND.n250 17.0005
R276 VGND.n260 VGND.n232 17.0005
R277 VGND.n260 VGND.n228 17.0005
R278 VGND.n260 VGND.n226 17.0005
R279 VGND.n260 VGND.n253 17.0005
R280 VGND.n493 VGND.n1 17.0005
R281 VGND.n494 VGND.n493 17.0005
R282 VGND.n489 VGND.n18 17.0005
R283 VGND.n489 VGND.n14 17.0005
R284 VGND.n489 VGND.n29 17.0005
R285 VGND.n489 VGND.n13 17.0005
R286 VGND.n489 VGND.n11 17.0005
R287 VGND.n489 VGND.n31 17.0005
R288 VGND.n484 VGND.n483 17.0005
R289 VGND.n483 VGND.n56 17.0005
R290 VGND.n483 VGND.n41 17.0005
R291 VGND.n483 VGND.n58 17.0005
R292 VGND.n483 VGND.n482 17.0005
R293 VGND.n288 VGND.n287 16.9935
R294 VGND.n270 VGND.n269 16.2915
R295 VGND.n269 VGND.n206 16.2014
R296 VGND.n474 VGND.n67 15.6652
R297 VGND.n284 VGND.n283 15.5838
R298 VGND.n396 VGND.n66 15.4962
R299 VGND.n297 VGND.n296 15.4044
R300 VGND.n479 VGND.n62 15.3111
R301 VGND.n206 VGND.n205 15.2207
R302 VGND.n271 VGND.n270 15.2126
R303 VGND.n351 VGND.n350 14.8829
R304 VGND.n209 VGND.n208 14.853
R305 VGND.n348 VGND.n347 14.853
R306 VGND.n294 VGND.n293 14.6742
R307 VGND.n296 VGND.n295 14.2225
R308 VGND.n477 VGND.n64 14.1685
R309 VGND.n285 VGND.n284 12.3693
R310 VGND.n496 VGND.n495 11.5981
R311 VGND.n410 VGND.n409 11.5903
R312 VGND.n451 VGND.n68 11.5621
R313 VGND.n278 VGND.n277 11.5336
R314 VGND.n75 VGND.n74 11.0666
R315 VGND.n469 VGND.n468 10.3577
R316 VGND.n198 VGND.n197 10.3577
R317 VGND.n377 VGND.n60 9.85117
R318 VGND.n195 VGND.n161 9.69267
R319 VGND.n439 VGND.n434 9.0005
R320 VGND.n434 VGND.n427 9.0005
R321 VGND.n439 VGND.n438 9.0005
R322 VGND.n438 VGND.n427 9.0005
R323 VGND.n439 VGND.n433 9.0005
R324 VGND.n440 VGND.n429 9.0005
R325 VGND.n440 VGND.n427 9.0005
R326 VGND.n440 VGND.n439 9.0005
R327 VGND.n445 VGND.n442 9.0005
R328 VGND.n442 VGND.n425 9.0005
R329 VGND.n445 VGND.n444 9.0005
R330 VGND.n444 VGND.n425 9.0005
R331 VGND.n445 VGND.n441 9.0005
R332 VGND.n447 VGND.n446 9.0005
R333 VGND.n446 VGND.n425 9.0005
R334 VGND.n446 VGND.n445 9.0005
R335 VGND.n446 uio_oe[7] 8.8478
R336 VGND.n44 VGND.t92 8.74885
R337 VGND.n26 VGND.t1 8.74885
R338 VGND.n247 VGND.t29 8.74885
R339 VGND.n239 VGND.n237 8.501
R340 VGND.n239 VGND.n238 8.501
R341 VGND.n492 VGND.n491 8.501
R342 VGND.n491 VGND.n6 8.501
R343 VGND.n52 VGND.n50 8.501
R344 VGND.n52 VGND.n51 8.501
R345 VGND.n264 VGND.n220 8.47111
R346 VGND.n263 VGND.n221 8.47111
R347 VGND.n262 VGND.n222 8.47111
R348 VGND.n260 VGND.n243 8.47111
R349 VGND.n260 VGND.n245 8.47111
R350 VGND.n260 VGND.n249 8.47111
R351 VGND.n260 VGND.n230 8.47111
R352 VGND.n260 VGND.n227 8.47111
R353 VGND.n260 VGND.n255 8.47111
R354 VGND.n4 VGND.n2 8.47111
R355 VGND.n17 VGND.n7 8.47111
R356 VGND.n489 VGND.n22 8.47111
R357 VGND.n489 VGND.n24 8.47111
R358 VGND.n489 VGND.n28 8.47111
R359 VGND.n489 VGND.n33 8.47111
R360 VGND.n487 VGND.n37 8.47111
R361 VGND.n486 VGND.n38 8.47111
R362 VGND.n485 VGND.n39 8.47111
R363 VGND.n483 VGND.n46 8.47111
R364 VGND.n483 VGND.n45 8.47111
R365 VGND.n483 VGND.n42 8.47111
R366 VGND.n273 VGND.n156 8.0799
R367 VGND.n464 VGND.n463 7.52168
R368 VGND.n464 VGND.n76 7.47272
R369 VGND.n281 VGND.n153 6.68645
R370 VGND.n398 VGND.n395 6.63864
R371 VGND.n467 VGND.n466 6.53659
R372 VGND.n163 VGND.n162 6.32858
R373 VGND.n192 VGND.n191 6.07977
R374 VGND.n196 VGND.n156 6.05718
R375 VGND.n273 VGND.n272 5.9638
R376 VGND.n240 VGND.n239 5.66778
R377 VGND.n491 VGND.n490 5.66778
R378 VGND.n52 VGND.n49 5.66778
R379 VGND.n239 VGND.n211 5.66767
R380 VGND.n491 VGND.n3 5.66767
R381 VGND.n52 VGND.n8 5.66767
R382 VGND.n260 VGND.n241 5.61485
R383 VGND.n260 VGND.n252 5.61485
R384 VGND.n489 VGND.n20 5.61485
R385 VGND.n489 VGND.n30 5.61485
R386 VGND.n483 VGND.n48 5.61485
R387 VGND.n291 VGND.n273 5.51412
R388 VGND.n433 VGND 5.4103
R389 VGND.n292 VGND.n291 4.6955
R390 VGND.n437 VGND.n436 4.49573
R391 VGND.n436 VGND.n428 4.49573
R392 VGND.n443 VGND.n400 4.49573
R393 VGND.n426 VGND.n400 4.49573
R394 VGND.n435 VGND.n429 4.49573
R395 VGND.n447 VGND.n403 4.49573
R396 VGND.n433 VGND.n432 4.4949
R397 VGND.n441 VGND.n402 4.4949
R398 VGND.n290 VGND.n289 4.09378
R399 VGND.n276 VGND.n274 3.42765
R400 VGND.n266 VGND.n216 3.38768
R401 VGND.n282 VGND.n281 3.27628
R402 VGND.n299 VGND.n298 2.85446
R403 VGND.n326 VGND.n125 2.31911
R404 VGND.n125 VGND 2.31911
R405 VGND.n78 VGND.n77 2.27849
R406 VGND.n449 VGND.n400 2.2505
R407 VGND.n448 VGND.n447 2.2505
R408 VGND.n436 VGND.n86 2.2505
R409 VGND.n430 VGND.n429 2.2505
R410 VGND.n266 VGND.n265 1.97699
R411 VGND.n260 VGND.n259 1.97699
R412 VGND.n489 VGND.n488 1.97699
R413 VGND.n311 VGND.n141 1.86972
R414 VGND.n453 VGND.n452 1.81263
R415 VGND.n346 VGND.n345 1.47805
R416 VGND.n345 VGND.n344 1.4745
R417 VGND.n399 VGND.n87 1.41597
R418 VGND.n441 VGND.n440 1.40696
R419 VGND.n260 VGND.n256 1.21402
R420 VGND.n489 VGND.n34 1.21402
R421 VGND.n266 VGND.n217 1.21402
R422 VGND.n281 VGND.n274 1.18201
R423 VGND.n448 VGND.n401 1.1463
R424 VGND.n431 VGND.n430 1.1463
R425 VGND.n398 VGND.n397 1.13055
R426 VGND.n89 VGND.n88 1.1093
R427 VGND.n266 VGND.n212 1.04263
R428 VGND.n260 VGND.n246 1.04263
R429 VGND.n260 VGND.n231 1.04263
R430 VGND.n260 VGND.n224 1.04263
R431 VGND.n489 VGND.n25 1.04263
R432 VGND.n489 VGND.n12 1.04263
R433 VGND.n489 VGND.n9 1.04263
R434 VGND.n483 VGND.n43 1.04263
R435 VGND.n260 VGND.n235 1.02715
R436 VGND.n260 VGND.n234 1.02715
R437 VGND.n489 VGND.n16 1.02715
R438 VGND.n489 VGND.n15 1.02715
R439 VGND.n483 VGND.n54 1.02715
R440 VGND.n483 VGND.n55 1.02715
R441 VGND.n328 VGND.n125 0.936079
R442 VGND.n207 VGND.n125 0.851167
R443 VGND.n353 VGND.n352 0.8068
R444 VGND.n379 VGND.n378 0.803036
R445 VGND.n399 VGND.n398 0.610292
R446 VGND.n383 VGND.n382 0.598489
R447 VGND.n311 VGND.n310 0.597922
R448 VGND.n265 VGND.n264 0.585769
R449 VGND.n488 VGND.n487 0.585769
R450 VGND.n259 VGND.n1 0.52548
R451 VGND.n450 VGND.n449 0.521717
R452 VGND.n465 VGND.n464 0.518224
R453 VGND.n265 VGND.n219 0.477006
R454 VGND.n259 VGND.n258 0.477006
R455 VGND.n488 VGND.n36 0.477006
R456 VGND.n345 VGND.n112 0.473781
R457 VGND.n163 VGND.n156 0.464095
R458 VGND.n455 VGND.n86 0.45348
R459 VGND.n341 VGND.n112 0.434656
R460 VGND.n384 VGND.n383 0.352948
R461 VGND.n310 VGND.n309 0.352948
R462 VGND.n341 VGND.n340 0.347746
R463 VGND.n164 VGND.n163 0.328048
R464 VGND.n291 VGND.n290 0.326045
R465 VGND.n404 uo_out[5] 0.32522
R466 VGND.n405 uo_out[6] 0.32522
R467 VGND.n406 uo_out[7] 0.32522
R468 VGND.n407 uio_out[0] 0.32522
R469 VGND.n412 uio_out[2] 0.32522
R470 VGND.n413 uio_out[3] 0.32522
R471 VGND.n414 uio_out[4] 0.32522
R472 VGND.n415 uio_out[5] 0.32522
R473 VGND.n416 uio_out[6] 0.32522
R474 VGND.n417 uio_out[7] 0.32522
R475 VGND.n418 uio_oe[0] 0.32522
R476 VGND.n419 uio_oe[1] 0.32522
R477 VGND.n420 uio_oe[2] 0.32522
R478 VGND.n421 uio_oe[3] 0.32522
R479 VGND.n422 uio_oe[4] 0.32522
R480 VGND.n423 uio_oe[5] 0.32522
R481 VGND.n424 uio_oe[6] 0.32522
R482 VGND.n340 VGND.n339 0.289181
R483 VGND.n496 VGND.n0 0.27022
R484 VGND.n385 VGND.n384 0.2683
R485 VGND.n309 VGND.n308 0.2683
R486 VGND.n189 VGND.n164 0.256021
R487 VGND.n344 VGND.n110 0.250193
R488 VGND.n453 VGND.n450 0.243514
R489 VGND.n339 VGND.n338 0.243383
R490 VGND.n264 VGND.n263 0.241078
R491 VGND.n263 VGND.n262 0.241078
R492 VGND.n17 VGND.n2 0.241078
R493 VGND.n487 VGND.n486 0.241078
R494 VGND.n486 VGND.n485 0.241078
R495 VGND.n411 VGND.n410 0.22226
R496 VGND.n386 VGND.n385 0.221084
R497 VGND.n308 VGND.n307 0.221084
R498 VGND.n338 VGND.n337 0.216589
R499 VGND.n219 VGND.n216 0.208
R500 VGND.n290 VGND.n274 0.201227
R501 VGND.n387 VGND.n386 0.193014
R502 VGND.n307 VGND.n306 0.193014
R503 VGND.n337 VGND.n336 0.189923
R504 VGND.n252 VGND 0.180825
R505 VGND.n30 VGND 0.180825
R506 VGND.n262 VGND.n261 0.180789
R507 VGND.n494 VGND.n2 0.180789
R508 VGND.n18 VGND.n17 0.180789
R509 VGND.n485 VGND.n484 0.180789
R510 VGND.n242 VGND.n241 0.177986
R511 VGND.n21 VGND.n20 0.177986
R512 VGND.n48 VGND.n47 0.177986
R513 VGND.n336 VGND.n335 0.177878
R514 VGND.n388 VGND.n387 0.172356
R515 VGND.n306 VGND.n305 0.172356
R516 VGND.n189 VGND.n188 0.165165
R517 VGND.n255 VGND.n254 0.163289
R518 VGND.n33 VGND.n32 0.163289
R519 VGND.n335 VGND.n334 0.161737
R520 VGND.n249 VGND.n248 0.159539
R521 VGND.n28 VGND.n27 0.159539
R522 VGND.n57 VGND.n42 0.159539
R523 VGND.n465 VGND.n73 0.158526
R524 VGND.n241 VGND.n223 0.158325
R525 VGND.n20 VGND.n19 0.158325
R526 VGND.n48 VGND.n40 0.158325
R527 VGND.n389 VGND.n388 0.155671
R528 VGND.n305 VGND.n304 0.155671
R529 VGND.n188 VGND.n187 0.152148
R530 VGND.n394 VGND.n393 0.150927
R531 VGND.n334 VGND.n333 0.149148
R532 VGND.n392 VGND.n90 0.149023
R533 VGND.n391 VGND.n91 0.147167
R534 VGND.n302 VGND.n150 0.147167
R535 VGND.n187 VGND.n186 0.145833
R536 VGND.n247 VGND.n245 0.145789
R537 VGND.n26 VGND.n24 0.145789
R538 VGND.n45 VGND.n44 0.145789
R539 VGND.n390 VGND.n92 0.144762
R540 VGND.n303 VGND.n149 0.144762
R541 VGND.n390 VGND.n389 0.143511
R542 VGND.n304 VGND.n303 0.143511
R543 VGND.n153 VGND.n152 0.143335
R544 VGND.n389 VGND.n93 0.14301
R545 VGND.n304 VGND.n148 0.14301
R546 VGND.n333 VGND.n332 0.142866
R547 VGND.n388 VGND.n94 0.1413
R548 VGND.n305 VGND.n147 0.1413
R549 VGND.n387 VGND.n95 0.13963
R550 VGND.n306 VGND.n146 0.13963
R551 VGND.n395 VGND.n89 0.139117
R552 VGND.n229 VGND.n227 0.138289
R553 VGND.n386 VGND.n96 0.138
R554 VGND.n307 VGND.n145 0.138
R555 VGND.n254 VGND.n252 0.137986
R556 VGND.n32 VGND.n30 0.137986
R557 VGND.n186 VGND.n185 0.136464
R558 VGND.n385 VGND.n97 0.136407
R559 VGND.n308 VGND.n144 0.136407
R560 VGND.n460 VGND.n459 0.134991
R561 VGND.n384 VGND.n98 0.134851
R562 VGND.n309 VGND.n143 0.134851
R563 VGND.n391 VGND.n390 0.134721
R564 VGND.n303 VGND.n302 0.134721
R565 VGND.n332 VGND.n331 0.133592
R566 VGND.n383 VGND.n99 0.13333
R567 VGND.n310 VGND.n142 0.13333
R568 VGND.n185 VGND.n184 0.131588
R569 VGND.n244 VGND.n243 0.130789
R570 VGND.n23 VGND.n22 0.130789
R571 VGND.n331 VGND.n330 0.127631
R572 VGND.n354 VGND.n109 0.127631
R573 VGND.n392 VGND.n391 0.127467
R574 VGND.n302 VGND.n301 0.127467
R575 VGND.n184 VGND.n183 0.126098
R576 VGND.n330 VGND.n329 0.123294
R577 VGND.n243 VGND.n242 0.123289
R578 VGND.n22 VGND.n21 0.123289
R579 VGND.n47 VGND.n46 0.123289
R580 VGND.n358 VGND.n109 0.122221
R581 VGND.n353 VGND.n110 0.122211
R582 VGND.n183 VGND.n182 0.121629
R583 VGND.n393 VGND.n392 0.121573
R584 VGND.n301 VGND.n300 0.121573
R585 VGND VGND.n230 0.120789
R586 VGND VGND.n227 0.120789
R587 VGND.n409 VGND.n46 0.120789
R588 VGND.n395 VGND.n394 0.119995
R589 VGND.n177 VGND.n176 0.119457
R590 VGND.n182 VGND.n181 0.118673
R591 VGND.n359 VGND.n358 0.117844
R592 VGND.n177 VGND.n73 0.117211
R593 VGND.n181 VGND.n180 0.114913
R594 VGND.n360 VGND.n359 0.114675
R595 VGND.n180 VGND.n179 0.113743
R596 VGND.n343 VGND.n112 0.112734
R597 VGND.n342 VGND.n341 0.112578
R598 VGND.n258 VGND.n255 0.112039
R599 VGND.n36 VGND.n33 0.112039
R600 VGND.n340 VGND.n113 0.111718
R601 VGND.n339 VGND.n114 0.111507
R602 VGND.n325 VGND.n324 0.111202
R603 VGND.n360 VGND.n107 0.111202
R604 VGND.n301 VGND.n151 0.11115
R605 VGND.n245 VGND.n244 0.110789
R606 VGND.n24 VGND.n23 0.110789
R607 VGND.n408 VGND.n45 0.110789
R608 VGND.n179 VGND.n178 0.110741
R609 VGND.n338 VGND.n115 0.110644
R610 VGND.n178 VGND.n177 0.110231
R611 VGND.n337 VGND.n116 0.110139
R612 VGND.n324 VGND.n323 0.110119
R613 VGND.n336 VGND.n117 0.109632
R614 VGND.n190 VGND.n189 0.109257
R615 VGND.n364 VGND.n107 0.109256
R616 VGND.n335 VGND.n118 0.109053
R617 VGND.n188 VGND.n165 0.10874
R618 VGND.n334 VGND.n119 0.10854
R619 VGND.n187 VGND.n166 0.108513
R620 VGND.n186 VGND.n167 0.108352
R621 VGND.n185 VGND.n168 0.108122
R622 VGND.n333 VGND.n120 0.108023
R623 VGND.n332 VGND.n121 0.107796
R624 VGND.n183 VGND.n170 0.107722
R625 VGND.n184 VGND.n169 0.107592
R626 VGND.n182 VGND.n171 0.107552
R627 VGND.n180 VGND.n173 0.10751
R628 VGND.n331 VGND.n122 0.107273
R629 VGND.n355 VGND.n354 0.107273
R630 VGND.n323 VGND.n322 0.107182
R631 VGND.n178 VGND.n175 0.107092
R632 VGND.n330 VGND.n123 0.107042
R633 VGND.n356 VGND.n109 0.107042
R634 VGND.n181 VGND.n172 0.10701
R635 VGND.n179 VGND.n174 0.106962
R636 VGND.n329 VGND.n124 0.10687
R637 VGND.n358 VGND.n357 0.10687
R638 VGND.n327 VGND.n126 0.106635
R639 VGND.n359 VGND.n108 0.106635
R640 VGND.n381 VGND.n101 0.106426
R641 VGND.n313 VGND.n139 0.106426
R642 VGND.n365 VGND.n364 0.106367
R643 VGND.n325 VGND.n127 0.1061
R644 VGND.n361 VGND.n360 0.1061
R645 VGND.n323 VGND.n129 0.10604
R646 VGND.n364 VGND.n363 0.10604
R647 VGND.n321 VGND.n131 0.105977
R648 VGND.n367 VGND.n366 0.105977
R649 VGND.n316 VGND.n136 0.105973
R650 VGND.n374 VGND.n103 0.105973
R651 VGND.n324 VGND.n128 0.10592
R652 VGND.n362 VGND.n107 0.10592
R653 VGND.n380 VGND.n102 0.105907
R654 VGND.n314 VGND.n138 0.105907
R655 VGND.n317 VGND.n135 0.105848
R656 VGND.n373 VGND.n372 0.105848
R657 VGND.n315 VGND.n137 0.10578
R658 VGND.n376 VGND.n375 0.10578
R659 VGND.n320 VGND.n132 0.105731
R660 VGND.n368 VGND.n105 0.105731
R661 VGND.n322 VGND.n321 0.105665
R662 VGND.n318 VGND.n134 0.105663
R663 VGND.n371 VGND.n104 0.105663
R664 VGND.n319 VGND.n133 0.105542
R665 VGND.n370 VGND.n369 0.105542
R666 VGND.n322 VGND.n130 0.105493
R667 VGND.n365 VGND.n106 0.105493
R668 VGND.n366 VGND.n365 0.104886
R669 VGND.n299 VGND.n153 0.104495
R670 VGND.n321 VGND.n320 0.104166
R671 VGND.n366 VGND.n105 0.104166
R672 VGND.n410 uio_out[1] 0.10346
R673 VGND.n230 VGND.n229 0.103289
R674 VGND.n319 VGND.n318 0.102551
R675 VGND.n320 VGND.n319 0.102053
R676 VGND.n370 VGND.n105 0.102053
R677 VGND.n326 VGND.n325 0.101891
R678 VGND.n371 VGND.n370 0.101858
R679 VGND.n318 VGND.n317 0.101493
R680 VGND.n372 VGND.n371 0.101493
R681 VGND.n317 VGND.n316 0.100967
R682 VGND.n372 VGND.n103 0.100967
R683 VGND.n314 VGND.n313 0.100958
R684 VGND.n315 VGND.n314 0.100445
R685 VGND.n381 VGND.n380 0.100376
R686 VGND.n316 VGND.n315 0.100187
R687 VGND.n376 VGND.n103 0.100187
R688 VGND.n73 VGND.n72 0.0973571
R689 VGND.n249 VGND.n247 0.095789
R690 VGND.n28 VGND.n26 0.095789
R691 VGND.n44 VGND.n42 0.095789
R692 VGND.n459 VGND.n458 0.0954338
R693 VGND.n454 VGND.n85 0.0928432
R694 VGND.n329 VGND.n328 0.0895217
R695 VGND.n463 VGND.n462 0.0873393
R696 VGND.n207 VGND 0.0854123
R697 VGND.n261 VGND.n223 0.083
R698 VGND.n19 VGND.n18 0.083
R699 VGND.n484 VGND.n40 0.083
R700 VGND.n382 VGND.n100 0.0802603
R701 VGND.n312 VGND.n140 0.0802603
R702 VGND.n101 VGND.n100 0.0782828
R703 VGND.n140 VGND.n139 0.0782828
R704 VGND.n495 VGND.n494 0.078
R705 VGND.n394 VGND.n90 0.0779701
R706 VGND.n380 VGND.n379 0.0771258
R707 VGND.n354 VGND.n353 0.0762778
R708 VGND.n458 VGND.n457 0.0754235
R709 VGND.n91 VGND.n90 0.0751329
R710 VGND.n454 VGND.n453 0.0739655
R711 VGND.n151 VGND.n150 0.0735315
R712 VGND.n92 VGND.n91 0.0731
R713 VGND.n150 VGND.n149 0.0731
R714 VGND.n462 VGND.n79 0.0724725
R715 VGND.n93 VGND.n92 0.0701066
R716 VGND.n149 VGND.n148 0.0701066
R717 VGND.n94 VGND.n93 0.067836
R718 VGND.n148 VGND.n147 0.067836
R719 VGND.n95 VGND.n94 0.06562
R720 VGND.n147 VGND.n146 0.06562
R721 VGND.n266 VGND.n213 0.0650946
R722 VGND.n260 VGND.n251 0.0650946
R723 VGND.n260 VGND.n225 0.0650946
R724 VGND.n489 VGND.n10 0.0650946
R725 VGND.n96 VGND.n95 0.0634565
R726 VGND.n146 VGND.n145 0.0634565
R727 VGND.n457 VGND.n456 0.0614573
R728 VGND.n292 VGND 0.061
R729 VGND.n272 VGND 0.061
R730 VGND.n397 VGND 0.061
R731 VGND.n77 VGND 0.061
R732 VGND.n76 VGND 0.061
R733 VGND.n467 VGND 0.061
R734 VGND.n192 VGND 0.061
R735 VGND.n162 VGND 0.061
R736 VGND.n452 VGND 0.061
R737 VGND.n87 VGND 0.061
R738 VGND.n88 VGND 0.061
R739 VGND.n97 VGND.n96 0.061
R740 VGND.n298 VGND 0.061
R741 VGND.n282 VGND 0.061
R742 VGND.n276 VGND 0.061
R743 VGND.n145 VGND.n144 0.061
R744 VGND.n141 VGND 0.061
R745 VGND.n346 VGND 0.061
R746 VGND.n352 VGND 0.061
R747 VGND.n378 VGND 0.061
R748 VGND.n196 VGND 0.061
R749 VGND.n289 VGND 0.061
R750 VGND.n81 VGND.n80 0.0607651
R751 VGND.n232 VGND 0.0605
R752 VGND VGND.n13 0.0605
R753 VGND.n58 VGND 0.0605
R754 VGND.n98 VGND.n97 0.0589402
R755 VGND.n144 VGND.n143 0.0589402
R756 VGND.n456 VGND.n455 0.0585315
R757 VGND.n300 VGND.n152 0.0568276
R758 VGND.n99 VGND.n98 0.0565916
R759 VGND.n143 VGND.n142 0.0565916
R760 uo_out[4] VGND.n496 0.0555
R761 VGND.n85 VGND.n84 0.0547113
R762 VGND.n100 VGND.n99 0.0546283
R763 VGND.n142 VGND.n140 0.0546283
R764 VGND.n460 VGND.n81 0.0545351
R765 VGND.n462 VGND.n461 0.0537058
R766 VGND.n382 VGND.n381 0.0505564
R767 VGND.n313 VGND.n312 0.0505564
R768 VGND.n102 VGND.n101 0.0497148
R769 VGND.n139 VGND.n138 0.0497148
R770 VGND.n84 VGND.n83 0.0483673
R771 VGND.n375 VGND.n102 0.0478846
R772 VGND.n138 VGND.n137 0.0478846
R773 VGND.n137 VGND.n136 0.04594
R774 VGND.n375 VGND.n374 0.04594
R775 VGND.n136 VGND.n135 0.0440235
R776 VGND.n374 VGND.n373 0.0440235
R777 VGND.n495 VGND.n1 0.043
R778 VGND.n450 VGND.n399 0.0425296
R779 VGND.n135 VGND.n134 0.0421344
R780 VGND.n373 VGND.n104 0.0421344
R781 VGND.n83 VGND.n82 0.0419304
R782 VGND.n176 VGND.n72 0.0411957
R783 VGND.n134 VGND.n133 0.0401312
R784 VGND.n369 VGND.n104 0.0401312
R785 VGND.n152 VGND.n151 0.0397586
R786 VGND.n393 VGND.n89 0.039235
R787 VGND.n133 VGND.n132 0.0386127
R788 VGND.n369 VGND.n368 0.0386127
R789 VGND.n132 VGND.n131 0.0365
R790 VGND.n368 VGND.n367 0.0365
R791 VGND.n466 VGND.n72 0.0356429
R792 VGND.n176 VGND.n175 0.0355141
R793 VGND.n131 VGND.n130 0.0351481
R794 VGND.n367 VGND.n106 0.0351481
R795 VGND.n175 VGND.n174 0.0337308
R796 VGND.n130 VGND.n129 0.0332724
R797 VGND.n363 VGND.n106 0.0332724
R798 VGND.n344 VGND.n343 0.032543
R799 VGND.n174 VGND.n173 0.0317753
R800 VGND.n129 VGND.n128 0.0313454
R801 VGND.n363 VGND.n362 0.0313454
R802 VGND.n355 VGND.n110 0.0307408
R803 VGND.n173 VGND.n172 0.0302379
R804 VGND.n128 VGND.n127 0.0299334
R805 VGND.n362 VGND.n361 0.0299334
R806 VGND.n328 VGND.n327 0.0298333
R807 VGND.n172 VGND.n171 0.0283213
R808 VGND.n127 VGND.n126 0.0279441
R809 VGND.n361 VGND.n108 0.0279441
R810 VGND.n80 VGND.n79 0.0273067
R811 VGND.n171 VGND.n170 0.0266297
R812 VGND.n126 VGND.n124 0.0263649
R813 VGND.n357 VGND.n108 0.0263649
R814 VGND.n170 VGND.n169 0.024961
R815 VGND.n447 VGND.n400 0.0249162
R816 VGND.n436 VGND.n429 0.0249162
R817 VGND.n124 VGND.n123 0.0247963
R818 VGND.n357 VGND.n356 0.0247963
R819 VGND.n169 VGND.n168 0.0233919
R820 VGND.n379 VGND.n376 0.02322
R821 VGND.n123 VGND.n122 0.0231622
R822 VGND.n356 VGND.n355 0.0231622
R823 VGND.n168 VGND.n167 0.0218333
R824 VGND.n248 VGND.n232 0.02175
R825 VGND.n27 VGND.n13 0.02175
R826 VGND.n58 VGND.n57 0.02175
R827 VGND.n449 VGND.n448 0.02162
R828 VGND.n430 VGND.n86 0.02162
R829 VGND.n122 VGND.n121 0.02162
R830 VGND.n466 VGND.n465 0.0212439
R831 VGND.n300 VGND.n299 0.0200345
R832 VGND.n167 VGND.n166 0.0199247
R833 VGND.n121 VGND.n120 0.0197957
R834 VGND.n166 VGND.n165 0.0186867
R835 VGND.n120 VGND.n119 0.0185662
R836 VGND.n461 VGND.n460 0.0170759
R837 VGND.n190 VGND.n165 0.0168721
R838 VGND.n119 VGND.n118 0.016764
R839 VGND.n0 uo_out[5] 0.0157601
R840 VGND.n404 uo_out[6] 0.0157601
R841 VGND.n405 uo_out[7] 0.0157601
R842 VGND.n406 uio_out[0] 0.0157601
R843 VGND.n407 uio_out[1] 0.0157601
R844 VGND.n411 uio_out[2] 0.0157601
R845 VGND.n412 uio_out[3] 0.0157601
R846 VGND.n413 uio_out[4] 0.0157601
R847 VGND.n414 uio_out[5] 0.0157601
R848 VGND.n415 uio_out[6] 0.0157601
R849 VGND.n416 uio_out[7] 0.0157601
R850 VGND.n417 uio_oe[0] 0.0157601
R851 VGND.n418 uio_oe[1] 0.0157601
R852 VGND.n419 uio_oe[2] 0.0157601
R853 VGND.n420 uio_oe[3] 0.0157601
R854 VGND.n421 uio_oe[4] 0.0157601
R855 VGND.n422 uio_oe[5] 0.0157601
R856 VGND.n423 uio_oe[6] 0.0157601
R857 VGND.n424 uio_oe[7] 0.0157601
R858 VGND.n79 VGND.n78 0.0153179
R859 VGND.n191 VGND.n190 0.0150695
R860 VGND.n118 VGND.n117 0.0149737
R861 VGND.n117 VGND.n116 0.0138158
R862 uo_out[5] VGND.n0 0.0137
R863 uo_out[6] VGND.n404 0.0137
R864 uo_out[7] VGND.n405 0.0137
R865 uio_out[0] VGND.n406 0.0137
R866 uio_out[1] VGND.n407 0.0137
R867 uio_out[2] VGND.n411 0.0137
R868 uio_out[3] VGND.n412 0.0137
R869 uio_out[4] VGND.n413 0.0137
R870 uio_out[5] VGND.n414 0.0137
R871 uio_out[6] VGND.n415 0.0137
R872 uio_out[7] VGND.n416 0.0137
R873 uio_oe[0] VGND.n417 0.0137
R874 uio_oe[1] VGND.n418 0.0137
R875 uio_oe[2] VGND.n419 0.0137
R876 uio_oe[3] VGND.n420 0.0137
R877 uio_oe[4] VGND.n421 0.0137
R878 uio_oe[5] VGND.n422 0.0137
R879 uio_oe[6] VGND.n423 0.0137
R880 uio_oe[7] VGND.n424 0.0137
R881 VGND.n327 VGND.n326 0.0132838
R882 VGND.n445 VGND.n401 0.0131992
R883 VGND.n439 VGND.n431 0.0131992
R884 VGND.n447 VGND.n402 0.0131916
R885 VGND.n432 VGND.n429 0.0131916
R886 VGND.n432 VGND.n427 0.0131916
R887 VGND.n425 VGND.n402 0.0131916
R888 VGND.n425 VGND.n401 0.0130858
R889 VGND.n431 VGND.n427 0.0130858
R890 VGND.n82 VGND.n81 0.0121797
R891 VGND.n116 VGND.n115 0.012041
R892 VGND.n446 VGND.n426 0.0115476
R893 VGND.n443 VGND.n441 0.0115476
R894 VGND.n440 VGND.n428 0.0115476
R895 VGND.n437 VGND.n433 0.0115476
R896 VGND.n434 VGND.n428 0.0115476
R897 VGND.n438 VGND.n437 0.0115476
R898 VGND.n442 VGND.n426 0.0115476
R899 VGND.n444 VGND.n443 0.0115476
R900 VGND.n444 VGND.n403 0.0115476
R901 VGND.n438 VGND.n435 0.0115476
R902 VGND.n435 VGND.n434 0.0115476
R903 VGND.n442 VGND.n403 0.0115476
R904 VGND.n115 VGND.n114 0.0105654
R905 VGND.n409 VGND.n408 0.0105
R906 VGND.n463 VGND.n78 0.00934499
R907 VGND.n455 VGND.n454 0.00920833
R908 VGND.n114 VGND.n113 0.00883987
R909 VGND.n459 VGND.n82 0.00874622
R910 VGND.n458 VGND.n83 0.0077971
R911 VGND.n342 VGND.n113 0.00737948
R912 VGND.n457 VGND.n84 0.00643951
R913 VGND.n343 VGND.n342 0.00594625
R914 VGND.n191 VGND.n164 0.00588981
R915 VGND.n461 VGND.n80 0.00446192
R916 VGND.n456 VGND.n85 0.00434654
R917 VGND.n312 VGND.n311 0.00206612
R918 VGND.n240 VGND.n222 0.00166667
R919 VGND.n490 VGND.n7 0.00166667
R920 VGND.n49 VGND.n39 0.00166667
R921 VGND.n260 VGND.n240 0.00133332
R922 VGND.n490 VGND.n489 0.00133332
R923 VGND.n483 VGND.n49 0.00133332
R924 VGND.n220 VGND.n211 0.001
R925 VGND.n237 VGND.n220 0.001
R926 VGND.n238 VGND.n221 0.001
R927 VGND.n493 VGND.n3 0.001
R928 VGND.n493 VGND.n492 0.001
R929 VGND.n6 VGND.n4 0.001
R930 VGND.n37 VGND.n8 0.001
R931 VGND.n50 VGND.n37 0.001
R932 VGND.n51 VGND.n38 0.001
R933 VGND.n266 VGND.n211 0.001
R934 VGND.n237 VGND.n221 0.001
R935 VGND.n238 VGND.n222 0.001
R936 VGND.n260 VGND.n3 0.001
R937 VGND.n492 VGND.n4 0.001
R938 VGND.n7 VGND.n6 0.001
R939 VGND.n489 VGND.n8 0.001
R940 VGND.n50 VGND.n38 0.001
R941 VGND.n51 VGND.n39 0.001
R942 uo_out[1].n3 uo_out[1].t2 15.0005
R943 uo_out[1] uo_out[1].n3 13.4668
R944 uo_out[1].n2 uo_out[1].n1 9.01747
R945 uo_out[1].n2 uo_out[1] 8.9065
R946 uo_out[1].n0 uo_out[1].t0 8.53421
R947 uo_out[1].n0 uo_out[1].t1 6.13626
R948 uo_out[1].n1 uo_out[1].n0 0.100612
R949 uo_out[1].n1 uo_out[1] 0.0585899
R950 uo_out[1].n3 uo_out[1] 0.04098
R951 uo_out[1] uo_out[1].n2 0.00678571
R952 VDPWR.n11 VDPWR.t48 34.1026
R953 VDPWR.n9 VDPWR.t14 34.1026
R954 VDPWR.n3 VDPWR.t10 34.1026
R955 VDPWR.n103 VDPWR.t29 34.1026
R956 VDPWR.n102 VDPWR.t67 34.1026
R957 VDPWR.n100 VDPWR.t56 34.1026
R958 VDPWR.n99 VDPWR.t46 34.1026
R959 VDPWR.n58 VDPWR.t6 34.1026
R960 VDPWR.n156 VDPWR.t21 34.1026
R961 VDPWR.n35 VDPWR.t72 34.1026
R962 VDPWR.n28 VDPWR.t42 34.1026
R963 VDPWR.n191 VDPWR.t58 34.1026
R964 VDPWR.n204 VDPWR.t36 34.1026
R965 VDPWR.n202 VDPWR.t50 34.1026
R966 VDPWR.n77 VDPWR.t17 34.1026
R967 VDPWR.n98 VDPWR.t44 34.1026
R968 VDPWR.n101 VDPWR.t64 34.1026
R969 VDPWR.n104 VDPWR.t33 34.1026
R970 VDPWR.n105 VDPWR.t4 34.1026
R971 VDPWR.n1 VDPWR.t62 34.1026
R972 VDPWR.n0 VDPWR.t8 34.1026
R973 VDPWR.n275 VDPWR.n214 19.7403
R974 VDPWR VDPWR.n11 18.2059
R975 VDPWR VDPWR.n9 18.2059
R976 VDPWR VDPWR.n3 18.2059
R977 VDPWR VDPWR.n103 18.2059
R978 VDPWR VDPWR.n102 18.2059
R979 VDPWR VDPWR.n100 18.2059
R980 VDPWR VDPWR.n99 18.2059
R981 VDPWR VDPWR.n58 18.2059
R982 VDPWR VDPWR.n156 18.2059
R983 VDPWR VDPWR.n35 18.2059
R984 VDPWR VDPWR.n28 18.2059
R985 VDPWR VDPWR.n191 18.2059
R986 VDPWR VDPWR.n204 18.2059
R987 VDPWR VDPWR.n202 18.2059
R988 VDPWR VDPWR.n77 18.2059
R989 VDPWR VDPWR.n98 18.2059
R990 VDPWR VDPWR.n101 18.2059
R991 VDPWR VDPWR.n104 18.2059
R992 VDPWR VDPWR.n105 18.2059
R993 VDPWR VDPWR.n1 18.2059
R994 VDPWR VDPWR.n0 18.2059
R995 VDPWR.n275 VDPWR.n274 18.0005
R996 VDPWR.n263 VDPWR.t66 17.378
R997 VDPWR.n248 VDPWR.t31 17.378
R998 VDPWR.n231 VDPWR.t35 17.378
R999 VDPWR.n264 VDPWR.t13 17.3693
R1000 VDPWR.n246 VDPWR.t27 17.3693
R1001 VDPWR.n230 VDPWR.t25 17.3693
R1002 VDPWR.n252 VDPWR.t3 17.1422
R1003 VDPWR.n11 VDPWR.t49 17.0233
R1004 VDPWR.n9 VDPWR.t15 17.0233
R1005 VDPWR.n3 VDPWR.t11 17.0233
R1006 VDPWR.n103 VDPWR.t30 17.0233
R1007 VDPWR.n102 VDPWR.t68 17.0233
R1008 VDPWR.n100 VDPWR.t57 17.0233
R1009 VDPWR.n99 VDPWR.t47 17.0233
R1010 VDPWR.n58 VDPWR.t7 17.0233
R1011 VDPWR.n156 VDPWR.t22 17.0233
R1012 VDPWR.n35 VDPWR.t73 17.0233
R1013 VDPWR.n28 VDPWR.t43 17.0233
R1014 VDPWR.n191 VDPWR.t59 17.0233
R1015 VDPWR.n204 VDPWR.t37 17.0233
R1016 VDPWR.n202 VDPWR.t51 17.0233
R1017 VDPWR.n77 VDPWR.t18 17.0233
R1018 VDPWR.n98 VDPWR.t45 17.0233
R1019 VDPWR.n101 VDPWR.t65 17.0233
R1020 VDPWR.n104 VDPWR.t34 17.0233
R1021 VDPWR.n105 VDPWR.t5 17.0233
R1022 VDPWR.n1 VDPWR.t63 17.0233
R1023 VDPWR.n0 VDPWR.t9 17.0233
R1024 VDPWR.n271 VDPWR.n229 17.0005
R1025 VDPWR.n272 VDPWR.n271 17.0005
R1026 VDPWR.n263 VDPWR.t16 17.0005
R1027 VDPWR.n248 VDPWR.t23 17.0005
R1028 VDPWR.n266 VDPWR.n250 17.0005
R1029 VDPWR.n266 VDPWR.n253 17.0005
R1030 VDPWR.n266 VDPWR.n254 17.0005
R1031 VDPWR.n266 VDPWR.n241 17.0005
R1032 VDPWR.n231 VDPWR.t28 17.0005
R1033 VDPWR.n271 VDPWR.n215 17.0005
R1034 VDPWR.n271 VDPWR.n222 17.0005
R1035 VDPWR.n271 VDPWR.n235 17.0005
R1036 VDPWR.n267 VDPWR.n266 17.0005
R1037 VDPWR.n276 VDPWR.n275 12.4694
R1038 VDPWR.n212 VDPWR.n211 9.2117
R1039 VDPWR.n208 VDPWR.n194 9.18823
R1040 VDPWR.n212 VDPWR.n22 9.18823
R1041 VDPWR.n212 VDPWR.n21 9.05079
R1042 VDPWR.n209 VDPWR.n208 9.0005
R1043 VDPWR.n210 VDPWR.n22 9.0005
R1044 VDPWR.n209 VDPWR.n25 9.0005
R1045 VDPWR.n210 VDPWR.n21 9.0005
R1046 VDPWR.n209 VDPWR.n23 9.0005
R1047 VDPWR.n211 VDPWR.n210 9.0005
R1048 VDPWR.n199 VDPWR.n198 9.0005
R1049 VDPWR.n196 VDPWR.n15 9.0005
R1050 VDPWR.n280 VDPWR.n17 9.0005
R1051 VDPWR.n261 VDPWR.t54 8.80285
R1052 VDPWR.n237 VDPWR.t75 8.80285
R1053 VDPWR.n225 VDPWR.t40 8.80285
R1054 VDPWR.t0 VDPWR.n242 8.501
R1055 VDPWR.n266 VDPWR.n258 8.47111
R1056 VDPWR.n266 VDPWR.n260 8.47111
R1057 VDPWR.n271 VDPWR.n226 8.47111
R1058 VDPWR.n271 VDPWR.n219 8.47111
R1059 VDPWR.n271 VDPWR.n217 8.47111
R1060 VDPWR.n269 VDPWR.n238 8.47111
R1061 VDPWR.n268 VDPWR.n239 8.47111
R1062 VDPWR.n259 VDPWR.t52 6.07323
R1063 VDPWR.n218 VDPWR.t74 6.07323
R1064 VDPWR.n224 VDPWR.t38 6.07323
R1065 VDPWR.n107 VDPWR.n106 6.01045
R1066 VDPWR.n228 VDPWR.t61 5.98925
R1067 VDPWR.n216 VDPWR.t60 5.98882
R1068 VDPWR.n257 VDPWR.t20 5.98882
R1069 VDPWR.n255 VDPWR.t19 5.98882
R1070 VDPWR.n220 VDPWR.t1 5.98882
R1071 VDPWR.n234 VDPWR.t2 5.98882
R1072 VDPWR.n109 VDPWR.n108 5.98145
R1073 VDPWR.n10 VDPWR 5.96901
R1074 VDPWR.n192 VDPWR.n190 5.84778
R1075 VDPWR.n271 VDPWR.n227 5.61485
R1076 VDPWR.n266 VDPWR.n251 5.61485
R1077 VDPWR.n266 VDPWR.n256 5.61485
R1078 VDPWR.n271 VDPWR.n221 5.61485
R1079 VDPWR.n271 VDPWR.n270 5.61485
R1080 VDPWR.n277 VDPWR 5.2541
R1081 VDPWR.n112 VDPWR.n111 5.21746
R1082 VDPWR.n4 VDPWR 4.89941
R1083 VDPWR.n284 VDPWR 4.6152
R1084 VDPWR.n194 VDPWR.n193 4.53071
R1085 VDPWR.n207 VDPWR.n26 4.51901
R1086 VDPWR.n206 VDPWR.n20 4.50989
R1087 VDPWR VDPWR.n295 4.13588
R1088 VDPWR.n2 VDPWR 3.92388
R1089 VDPWR.n107 VDPWR 3.88095
R1090 VDPWR.n106 VDPWR 3.84419
R1091 VDPWR.n203 VDPWR 3.78722
R1092 VDPWR.n108 VDPWR 3.41222
R1093 VDPWR.n271 VDPWR.n233 3.30723
R1094 VDPWR.n266 VDPWR.n247 3.30688
R1095 VDPWR.n205 VDPWR 3.28289
R1096 VDPWR.n198 VDPWR.n197 3.0005
R1097 VDPWR.n15 VDPWR.n13 3.0005
R1098 VDPWR.n281 VDPWR.n280 3.0005
R1099 VDPWR.n192 VDPWR 2.98934
R1100 VDPWR.n266 VDPWR.n265 2.72512
R1101 VDPWR.n284 VDPWR.n283 2.5318
R1102 VDPWR.n29 VDPWR 2.53128
R1103 VDPWR.n155 VDPWR.n57 2.46388
R1104 VDPWR.n109 VDPWR 2.33518
R1105 VDPWR.n266 VDPWR.n245 2.29781
R1106 VDPWR.n194 VDPWR.n24 2.27162
R1107 VDPWR.n195 VDPWR.n16 2.26628
R1108 VDPWR.n213 VDPWR.n212 2.2505
R1109 VDPWR.n209 VDPWR.n24 2.2505
R1110 VDPWR.n210 VDPWR.n19 2.2505
R1111 VDPWR.n278 VDPWR.n16 2.2505
R1112 VDPWR.n280 VDPWR.n279 2.2505
R1113 VDPWR.n244 VDPWR 2.0605
R1114 VDPWR.n36 VDPWR 1.94477
R1115 VDPWR.n277 VDPWR.n276 1.89976
R1116 VDPWR.n110 VDPWR 1.74056
R1117 VDPWR.n112 VDPWR 1.53994
R1118 VDPWR.n240 VDPWR 1.53643
R1119 VDPWR.n278 VDPWR.n277 1.47736
R1120 VDPWR.n276 VDPWR.n213 1.46416
R1121 VDPWR.n111 VDPWR 1.39911
R1122 VDPWR.n157 VDPWR 1.30374
R1123 VDPWR.n114 VDPWR 1.19117
R1124 VDPWR.n279 VDPWR.n18 1.14638
R1125 VDPWR.n113 VDPWR.n112 0.923201
R1126 VDPWR.n135 VDPWR 0.895684
R1127 VDPWR.n154 VDPWR 0.886
R1128 VDPWR.n225 VDPWR.n223 0.854038
R1129 VDPWR.n262 VDPWR.n261 0.851125
R1130 VDPWR.n264 VDPWR.n262 0.805789
R1131 VDPWR.n230 VDPWR.n223 0.803932
R1132 VDPWR.n271 VDPWR.n223 0.802654
R1133 VDPWR.n266 VDPWR.n262 0.800901
R1134 VDPWR.n295 VDPWR.n294 0.762687
R1135 VDPWR.n273 VDPWR 0.543
R1136 VDPWR.n185 VDPWR.n27 0.531002
R1137 VDPWR.n169 VDPWR.n168 0.507992
R1138 VDPWR.n84 VDPWR.n83 0.507992
R1139 VDPWR.n265 VDPWR.n263 0.410237
R1140 VDPWR.n110 VDPWR.n109 0.409089
R1141 VDPWR.t0 VDPWR.n236 0.40574
R1142 VDPWR.n245 VDPWR.n244 0.392462
R1143 VDPWR.n265 VDPWR.n264 0.389189
R1144 VDPWR.n246 VDPWR.n245 0.373903
R1145 VDPWR.n106 VDPWR.n2 0.363276
R1146 VDPWR.n205 VDPWR.n203 0.348974
R1147 VDPWR.n243 VDPWR.t0 0.341
R1148 VDPWR.n233 VDPWR.n230 0.336433
R1149 VDPWR.n247 VDPWR.n246 0.335808
R1150 VDPWR.n111 VDPWR.n110 0.332665
R1151 VDPWR.n249 VDPWR.n247 0.332049
R1152 VDPWR.n233 VDPWR.n232 0.331445
R1153 VDPWR.n59 VDPWR.n57 0.330588
R1154 VDPWR.n108 VDPWR.n107 0.323555
R1155 VDPWR.n158 VDPWR.n155 0.313098
R1156 VDPWR.n206 VDPWR.n205 0.312824
R1157 VDPWR.n270 VDPWR.n269 0.300775
R1158 VDPWR.n295 VDPWR.n2 0.289257
R1159 VDPWR.n170 VDPWR.n169 0.2887
R1160 VDPWR.n85 VDPWR.n84 0.2887
R1161 VDPWR.n60 VDPWR.n59 0.280623
R1162 VDPWR.n184 VDPWR.n30 0.251853
R1163 VDPWR.n183 VDPWR.n31 0.2469
R1164 VDPWR.n182 VDPWR.n32 0.24161
R1165 VDPWR.n115 VDPWR.n97 0.24161
R1166 VDPWR.n269 VDPWR.n268 0.241078
R1167 VDPWR.n61 VDPWR.n60 0.240286
R1168 VDPWR.n181 VDPWR.n33 0.237849
R1169 VDPWR.n116 VDPWR.n96 0.237849
R1170 VDPWR.n180 VDPWR.n34 0.234669
R1171 VDPWR.n117 VDPWR.n95 0.234669
R1172 VDPWR.n252 VDPWR.n251 0.234575
R1173 VDPWR.n179 VDPWR.n36 0.231561
R1174 VDPWR.n118 VDPWR.n94 0.231561
R1175 VDPWR.n189 VDPWR.n188 0.230306
R1176 VDPWR.n178 VDPWR.n37 0.226786
R1177 VDPWR.n119 VDPWR.n93 0.226786
R1178 VDPWR.n171 VDPWR.n170 0.225081
R1179 VDPWR.n86 VDPWR.n85 0.225081
R1180 VDPWR.n177 VDPWR.n38 0.22337
R1181 VDPWR.n120 VDPWR.n92 0.22337
R1182 VDPWR.n176 VDPWR.n39 0.219324
R1183 VDPWR.n121 VDPWR.n91 0.219324
R1184 VDPWR.n175 VDPWR.n40 0.217223
R1185 VDPWR.n122 VDPWR.n90 0.217223
R1186 VDPWR.n174 VDPWR.n41 0.213359
R1187 VDPWR.n123 VDPWR.n89 0.213359
R1188 VDPWR.n186 VDPWR.n185 0.212767
R1189 VDPWR.n211 VDPWR.n23 0.2117
R1190 VDPWR.n173 VDPWR.n42 0.211333
R1191 VDPWR.n124 VDPWR.n88 0.211333
R1192 VDPWR.n172 VDPWR.n43 0.208253
R1193 VDPWR.n125 VDPWR.n87 0.208253
R1194 VDPWR.n62 VDPWR.n61 0.204702
R1195 VDPWR.n171 VDPWR.n44 0.204642
R1196 VDPWR.n126 VDPWR.n86 0.204642
R1197 VDPWR.n170 VDPWR.n45 0.202722
R1198 VDPWR.n127 VDPWR.n85 0.202722
R1199 VDPWR.n190 VDPWR.n27 0.201278
R1200 VDPWR.n169 VDPWR.n46 0.19982
R1201 VDPWR.n128 VDPWR.n84 0.19982
R1202 VDPWR.n159 VDPWR.n158 0.193685
R1203 VDPWR.n63 VDPWR.n62 0.187779
R1204 VDPWR.n270 VDPWR.n237 0.185825
R1205 VDPWR.n268 VDPWR.n267 0.180789
R1206 VDPWR.n251 VDPWR 0.180486
R1207 VDPWR.n172 VDPWR.n171 0.177266
R1208 VDPWR.n87 VDPWR.n86 0.177266
R1209 VDPWR.n64 VDPWR.n63 0.175509
R1210 VDPWR.n167 VDPWR.n48 0.173049
R1211 VDPWR.n130 VDPWR.n82 0.173049
R1212 VDPWR.n166 VDPWR.n49 0.172207
R1213 VDPWR.n131 VDPWR.n81 0.172207
R1214 VDPWR.n258 VDPWR.n257 0.172039
R1215 VDPWR.n220 VDPWR.n219 0.172039
R1216 VDPWR.n165 VDPWR.n50 0.171374
R1217 VDPWR.n132 VDPWR.n80 0.171374
R1218 VDPWR.n164 VDPWR.n51 0.169731
R1219 VDPWR.n133 VDPWR.n79 0.169731
R1220 VDPWR.n163 VDPWR.n52 0.168921
R1221 VDPWR.n134 VDPWR.n78 0.168921
R1222 VDPWR.n201 VDPWR.n200 0.168402
R1223 VDPWR.n162 VDPWR.n53 0.167325
R1224 VDPWR.n135 VDPWR.n76 0.167325
R1225 VDPWR.n294 VDPWR.n293 0.166596
R1226 VDPWR.n161 VDPWR.n54 0.166538
R1227 VDPWR.n136 VDPWR.n75 0.166538
R1228 VDPWR.n160 VDPWR.n55 0.165758
R1229 VDPWR.n137 VDPWR.n74 0.165758
R1230 VDPWR.n113 VDPWR.n97 0.165337
R1231 VDPWR.n159 VDPWR.n56 0.164986
R1232 VDPWR.n138 VDPWR.n73 0.164986
R1233 VDPWR.n139 VDPWR.n72 0.164221
R1234 VDPWR.n140 VDPWR.n71 0.163463
R1235 VDPWR.n188 VDPWR.n187 0.162204
R1236 VDPWR.n142 VDPWR.n69 0.161968
R1237 VDPWR.n141 VDPWR.n70 0.161968
R1238 VDPWR.n144 VDPWR.n67 0.161231
R1239 VDPWR.n143 VDPWR.n68 0.161231
R1240 VDPWR.n147 VDPWR.n64 0.159776
R1241 VDPWR.n146 VDPWR.n65 0.159776
R1242 VDPWR.n145 VDPWR.n66 0.159776
R1243 VDPWR.n149 VDPWR.n62 0.159059
R1244 VDPWR.n148 VDPWR.n63 0.159059
R1245 VDPWR.n152 VDPWR.n59 0.158348
R1246 VDPWR.n151 VDPWR.n60 0.158348
R1247 VDPWR.n150 VDPWR.n61 0.158348
R1248 VDPWR.n65 VDPWR.n64 0.157911
R1249 VDPWR.n173 VDPWR.n172 0.157621
R1250 VDPWR.n88 VDPWR.n87 0.157621
R1251 VDPWR.n153 VDPWR.n57 0.154546
R1252 VDPWR.n168 VDPWR.n47 0.15242
R1253 VDPWR.n129 VDPWR.n83 0.15242
R1254 VDPWR.n286 VDPWR.n285 0.152188
R1255 VDPWR.n66 VDPWR.n65 0.147308
R1256 VDPWR.n207 VDPWR.n22 0.147167
R1257 VDPWR.n67 VDPWR.n66 0.14126
R1258 VDPWR.n174 VDPWR.n173 0.141098
R1259 VDPWR.n89 VDPWR.n88 0.141098
R1260 VDPWR.n260 VDPWR.n259 0.140789
R1261 VDPWR.n218 VDPWR.n217 0.140789
R1262 VDPWR.n226 VDPWR.n224 0.140789
R1263 VDPWR.n294 VDPWR.n4 0.137615
R1264 VDPWR.n249 VDPWR.n248 0.136382
R1265 VDPWR.n232 VDPWR.n231 0.136382
R1266 VDPWR.n291 VDPWR.n5 0.135022
R1267 VDPWR.n68 VDPWR.n67 0.133682
R1268 VDPWR.n227 VDPWR.n216 0.129236
R1269 VDPWR.n257 VDPWR.n256 0.129236
R1270 VDPWR.n221 VDPWR.n220 0.129236
R1271 VDPWR.n228 VDPWR.n227 0.128325
R1272 VDPWR.n256 VDPWR.n255 0.128325
R1273 VDPWR.n234 VDPWR.n221 0.128325
R1274 VDPWR.n69 VDPWR.n68 0.127233
R1275 VDPWR.n186 VDPWR.n30 0.1269
R1276 VDPWR.n175 VDPWR.n174 0.126475
R1277 VDPWR.n90 VDPWR.n89 0.126475
R1278 VDPWR.n70 VDPWR.n69 0.123269
R1279 VDPWR.n71 VDPWR.n70 0.121562
R1280 VDPWR.n193 VDPWR.n23 0.1171
R1281 VDPWR.n72 VDPWR.n71 0.116891
R1282 VDPWR.n176 VDPWR.n175 0.116337
R1283 VDPWR.n91 VDPWR.n90 0.116337
R1284 VDPWR.n261 VDPWR.n260 0.115789
R1285 VDPWR.n237 VDPWR.n217 0.115789
R1286 VDPWR.n226 VDPWR.n225 0.115789
R1287 VDPWR.n73 VDPWR.n72 0.114401
R1288 VDPWR.n229 VDPWR.n228 0.113
R1289 VDPWR.n255 VDPWR.n254 0.113
R1290 VDPWR.n235 VDPWR.n234 0.113
R1291 VDPWR.n272 VDPWR.n216 0.11175
R1292 VDPWR.n160 VDPWR.n159 0.111106
R1293 VDPWR.n74 VDPWR.n73 0.111106
R1294 VDPWR.n161 VDPWR.n160 0.110556
R1295 VDPWR.n75 VDPWR.n74 0.110556
R1296 VDPWR.n162 VDPWR.n161 0.108981
R1297 VDPWR.n76 VDPWR.n75 0.108981
R1298 VDPWR.n78 VDPWR.n76 0.108669
R1299 VDPWR.n79 VDPWR.n78 0.108583
R1300 VDPWR.n177 VDPWR.n176 0.108277
R1301 VDPWR.n92 VDPWR.n91 0.108277
R1302 VDPWR.n80 VDPWR.n79 0.108072
R1303 VDPWR.n163 VDPWR.n162 0.107646
R1304 VDPWR.n164 VDPWR.n163 0.107594
R1305 VDPWR.n82 VDPWR.n81 0.107345
R1306 VDPWR.n166 VDPWR.n165 0.107234
R1307 VDPWR.n81 VDPWR.n80 0.107234
R1308 VDPWR.n165 VDPWR.n164 0.107115
R1309 VDPWR.n167 VDPWR.n166 0.106465
R1310 VDPWR.n178 VDPWR.n177 0.103826
R1311 VDPWR.n93 VDPWR.n92 0.103826
R1312 VDPWR.n259 VDPWR.n258 0.100789
R1313 VDPWR.n219 VDPWR.n218 0.100789
R1314 VDPWR.n179 VDPWR.n178 0.0994295
R1315 VDPWR.n94 VDPWR.n93 0.0994295
R1316 VDPWR.n180 VDPWR.n179 0.096586
R1317 VDPWR.n95 VDPWR.n94 0.096586
R1318 VDPWR.n288 VDPWR.n8 0.0942964
R1319 VDPWR.n181 VDPWR.n180 0.0929227
R1320 VDPWR.n96 VDPWR.n95 0.0929227
R1321 VDPWR.n182 VDPWR.n181 0.0912154
R1322 VDPWR.n97 VDPWR.n96 0.0912154
R1323 VDPWR.n6 VDPWR.n5 0.0893224
R1324 VDPWR.n183 VDPWR.n182 0.0884738
R1325 VDPWR.n274 VDPWR.n273 0.088
R1326 VDPWR.n184 VDPWR.n183 0.0871337
R1327 VDPWR.n185 VDPWR.n184 0.0864426
R1328 VDPWR.n31 VDPWR.n30 0.0816497
R1329 VDPWR.n187 VDPWR.n186 0.0787288
R1330 VDPWR.n32 VDPWR.n31 0.0781471
R1331 VDPWR.n115 VDPWR.n114 0.0781471
R1332 VDPWR.n292 VDPWR.n291 0.0761377
R1333 VDPWR.n33 VDPWR.n32 0.0757832
R1334 VDPWR.n116 VDPWR.n115 0.0757832
R1335 VDPWR.n34 VDPWR.n33 0.0734143
R1336 VDPWR.n117 VDPWR.n116 0.0734143
R1337 VDPWR.n291 VDPWR.n290 0.0722058
R1338 VDPWR.n240 VDPWR.n214 0.0717963
R1339 VDPWR.n287 VDPWR.n10 0.071653
R1340 VDPWR.n36 VDPWR.n34 0.071596
R1341 VDPWR.n118 VDPWR.n117 0.071596
R1342 VDPWR.n37 VDPWR.n36 0.0688352
R1343 VDPWR.n119 VDPWR.n118 0.0688352
R1344 VDPWR.n48 VDPWR.n47 0.0683607
R1345 VDPWR.n130 VDPWR.n129 0.0683607
R1346 VDPWR.n288 VDPWR.n287 0.0679195
R1347 VDPWR.n38 VDPWR.n37 0.0662582
R1348 VDPWR.n120 VDPWR.n119 0.0662582
R1349 VDPWR.n244 VDPWR.n241 0.0656852
R1350 VDPWR.n188 VDPWR.n27 0.0656852
R1351 VDPWR.n39 VDPWR.n38 0.0641087
R1352 VDPWR.n121 VDPWR.n120 0.0641087
R1353 VDPWR.n114 VDPWR.n113 0.0637952
R1354 VDPWR.n197 VDPWR.n12 0.0627642
R1355 VDPWR.n200 VDPWR.n199 0.0624718
R1356 VDPWR.n40 VDPWR.n39 0.0612059
R1357 VDPWR.n122 VDPWR.n121 0.0612059
R1358 VDPWR.n229 VDPWR 0.0605
R1359 VDPWR.n254 VDPWR 0.0605
R1360 VDPWR VDPWR.n253 0.0605
R1361 VDPWR VDPWR.n250 0.0605
R1362 VDPWR.n235 VDPWR 0.0605
R1363 VDPWR VDPWR.n222 0.0605
R1364 VDPWR.n41 VDPWR.n40 0.0599468
R1365 VDPWR.n123 VDPWR.n122 0.0599468
R1366 VDPWR.n289 VDPWR.n7 0.0577377
R1367 VDPWR.n42 VDPWR.n41 0.0571702
R1368 VDPWR.n124 VDPWR.n123 0.0571702
R1369 VDPWR.n43 VDPWR.n42 0.0555
R1370 VDPWR.n125 VDPWR.n124 0.0555
R1371 VDPWR.n44 VDPWR.n43 0.0535722
R1372 VDPWR.n126 VDPWR.n125 0.0535722
R1373 VDPWR.n285 VDPWR.n284 0.0532395
R1374 VDPWR.n292 VDPWR.n4 0.0528027
R1375 VDPWR.n293 VDPWR.n292 0.0522
R1376 VDPWR.n45 VDPWR.n44 0.0509772
R1377 VDPWR.n127 VDPWR.n126 0.0509772
R1378 VDPWR.n46 VDPWR.n45 0.0493889
R1379 VDPWR.n128 VDPWR.n127 0.0493889
R1380 VDPWR.n47 VDPWR.n46 0.04758
R1381 VDPWR.n129 VDPWR.n128 0.04758
R1382 VDPWR.n283 VDPWR.n12 0.0460752
R1383 VDPWR.n190 VDPWR.n189 0.045577
R1384 VDPWR.n168 VDPWR.n167 0.0448348
R1385 VDPWR.n83 VDPWR.n82 0.0448348
R1386 VDPWR.n49 VDPWR.n48 0.0427745
R1387 VDPWR.n131 VDPWR.n130 0.0427745
R1388 VDPWR.n287 VDPWR.n286 0.0419028
R1389 VDPWR.n208 VDPWR.n207 0.0415667
R1390 VDPWR.n200 VDPWR.n12 0.0413571
R1391 VDPWR.n289 VDPWR.n288 0.0410333
R1392 VDPWR.n283 VDPWR.n282 0.0408577
R1393 VDPWR.n50 VDPWR.n49 0.0408512
R1394 VDPWR.n132 VDPWR.n131 0.0408512
R1395 VDPWR.n224 VDPWR.n215 0.0405
R1396 VDPWR.n197 VDPWR.n13 0.0403491
R1397 VDPWR.n199 VDPWR.n196 0.040162
R1398 VDPWR.n196 VDPWR.n17 0.040162
R1399 VDPWR.n207 VDPWR.n21 0.0397857
R1400 VDPWR.n51 VDPWR.n50 0.0389466
R1401 VDPWR.n133 VDPWR.n132 0.0389466
R1402 VDPWR.n207 VDPWR.n206 0.0385976
R1403 VDPWR.n187 VDPWR.n29 0.0383925
R1404 VDPWR.n52 VDPWR.n51 0.0377308
R1405 VDPWR.n134 VDPWR.n133 0.0377308
R1406 VDPWR.n189 VDPWR.n29 0.0376329
R1407 VDPWR.n53 VDPWR.n52 0.0358684
R1408 VDPWR.n135 VDPWR.n134 0.0358684
R1409 VDPWR.n290 VDPWR.n289 0.0356133
R1410 VDPWR.n282 VDPWR.n13 0.0341226
R1411 VDPWR.n54 VDPWR.n53 0.0338649
R1412 VDPWR.n136 VDPWR.n135 0.0338649
R1413 VDPWR.n55 VDPWR.n54 0.0320472
R1414 VDPWR.n137 VDPWR.n136 0.0320472
R1415 VDPWR.n56 VDPWR.n55 0.0306596
R1416 VDPWR.n138 VDPWR.n137 0.0306596
R1417 VDPWR.n274 VDPWR.n215 0.0305
R1418 VDPWR.n157 VDPWR.n56 0.0288738
R1419 VDPWR.n139 VDPWR.n138 0.0288738
R1420 VDPWR.n193 VDPWR.n25 0.0282619
R1421 VDPWR.n140 VDPWR.n139 0.0271047
R1422 VDPWR.n250 VDPWR.n249 0.02675
R1423 VDPWR.n232 VDPWR.n222 0.02675
R1424 VDPWR.n141 VDPWR.n140 0.0257593
R1425 VDPWR.n267 VDPWR.n240 0.0255
R1426 VDPWR.n210 VDPWR.n209 0.0249162
R1427 VDPWR.n280 VDPWR.n15 0.0249162
R1428 VDPWR.n280 VDPWR.n16 0.0249162
R1429 VDPWR.n142 VDPWR.n141 0.0239128
R1430 VDPWR.n155 VDPWR.n154 0.02261
R1431 VDPWR.n203 VDPWR.n201 0.0225381
R1432 VDPWR.n143 VDPWR.n142 0.0222982
R1433 VDPWR.n24 VDPWR.n19 0.02162
R1434 VDPWR.n213 VDPWR.n19 0.02162
R1435 VDPWR.n279 VDPWR.n278 0.02162
R1436 VDPWR.n144 VDPWR.n143 0.0205913
R1437 VDPWR.n145 VDPWR.n144 0.018984
R1438 VDPWR.n286 VDPWR.n8 0.0188236
R1439 VDPWR.n158 VDPWR.n157 0.018557
R1440 VDPWR.n193 VDPWR.n192 0.0182408
R1441 VDPWR.n154 VDPWR.n153 0.0179271
R1442 VDPWR.n146 VDPWR.n145 0.0176222
R1443 VDPWR.n201 VDPWR.n195 0.0170391
R1444 VDPWR.n147 VDPWR.n146 0.0160294
R1445 VDPWR.n293 VDPWR.n5 0.015852
R1446 VDPWR.n8 VDPWR.n7 0.0156247
R1447 VDPWR.n285 VDPWR.n10 0.0149236
R1448 VDPWR.n7 VDPWR.n6 0.0148367
R1449 VDPWR.n148 VDPWR.n147 0.0140385
R1450 VDPWR.n198 VDPWR.n18 0.0138871
R1451 VDPWR.n18 VDPWR.n15 0.0133938
R1452 VDPWR.n194 VDPWR.n26 0.0132264
R1453 VDPWR.n212 VDPWR.n20 0.0132264
R1454 VDPWR.n149 VDPWR.n148 0.0131847
R1455 VDPWR.n209 VDPWR.n26 0.0131568
R1456 VDPWR.n210 VDPWR.n20 0.0131568
R1457 VDPWR.n207 VDPWR.n25 0.0115
R1458 VDPWR.n150 VDPWR.n149 0.0112027
R1459 VDPWR.n281 VDPWR.n14 0.0100472
R1460 VDPWR.n17 VDPWR.n14 0.0100023
R1461 VDPWR.n151 VDPWR.n150 0.00957623
R1462 VDPWR.n152 VDPWR.n151 0.00839238
R1463 VDPWR.n253 VDPWR.n252 0.00675
R1464 VDPWR.n282 VDPWR.n281 0.00672642
R1465 VDPWR.n241 VDPWR.n214 0.00661111
R1466 VDPWR.n153 VDPWR.n152 0.00641928
R1467 VDPWR.n195 VDPWR.n14 0.00463323
R1468 VDPWR.n273 VDPWR.n272 0.003
R1469 VDPWR.n238 VDPWR.n236 0.00197617
R1470 VDPWR.n290 VDPWR.n6 0.00108355
R1471 VDPWR.n271 VDPWR.n236 0.00102381
R1472 VDPWR.n243 VDPWR.n239 0.001
R1473 VDPWR.n242 VDPWR.n239 0.001
R1474 VDPWR.n266 VDPWR.n243 0.001
R1475 VDPWR.n242 VDPWR.n238 0.001
R1476 uo_out[2].n3 uo_out[2].t2 15.0005
R1477 uo_out[2] uo_out[2].n3 12.8496
R1478 uo_out[2].n2 uo_out[2] 12.5614
R1479 uo_out[2].n2 uo_out[2].n1 9.01936
R1480 uo_out[2].n0 uo_out[2].t0 8.53421
R1481 uo_out[2].n0 uo_out[2].t1 6.13626
R1482 uo_out[2].n1 uo_out[2].n0 0.0993764
R1483 uo_out[2].n1 uo_out[2] 0.0598258
R1484 uo_out[2] uo_out[2].n2 0.0388429
R1485 uo_out[2].n3 uo_out[2] 0.02525
R1486 uo_out[0].n4 uo_out[0].n3 33.1637
R1487 uo_out[0].n5 uo_out[0].t0 18.0455
R1488 uo_out[0] uo_out[0].t1 18.0125
R1489 uo_out[0].n1 uo_out[0].t3 15.0005
R1490 uo_out[0].n2 uo_out[0].n1 9.03505
R1491 uo_out[0].n3 uo_out[0].n2 6.7505
R1492 uo_out[0].n5 uo_out[0].n4 6.67645
R1493 uo_out[0].n4 uo_out[0].n0 4.90955
R1494 uo_out[0].n0 uo_out[0].t2 3.93974
R1495 uo_out[0].n3 uo_out[0] 1.35863
R1496 uo_out[0] uo_out[0].n5 0.0885
R1497 uo_out[0].n0 uo_out[0] 0.0446962
R1498 uo_out[0].n2 uo_out[0] 0.0401
R1499 uo_out[0].n1 uo_out[0] 0.02525
R1500 uo_out[3].n2 uo_out[3] 15.6957
R1501 uo_out[3].n2 uo_out[3].n1 9.0225
R1502 uo_out[3].n0 uo_out[3].t0 8.53421
R1503 uo_out[3].n0 uo_out[3].t1 6.13626
R1504 uo_out[3].n1 uo_out[3].n0 0.11668
R1505 uo_out[3].n1 uo_out[3] 0.0425225
R1506 uo_out[3] uo_out[3].n2 0.0357
C10 uo_out[0] VGND 11.2452f
C11 VDPWR VGND 0.10246p
.ends

