* NGSPICE file created from tt_um_oscillating_bones.ext - technology: ihp-sg13g2

.subckt tt_um_oscillating_bones ena clk rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] VGND VDPWR
X0 uo_out[1].t0 a_22205_61585# VGND.t119 VGND.t118 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X1 VDPWR.t52 a_16367_61578# freq_divider_0.sg13g2_dfrbp_2_0.D VDPWR.t2 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X2 VGND.t18 a_17996_61559# a_17075_61640# VGND.t37 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X3 VGND.t30 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_21132_61704# VGND.t29 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X4 a_16707_61717# a_16367_61578# VDPWR.t52 VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X5 a_17910_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t20 VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X6 a_20876_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t19 VDPWR.t2 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X7 ring_0/inverter_ring_0/skullfet_inverter_19.A ring_0/inverter_ring_0/skullfet_inverter_0.Y VDPWR.t44 VDPWR.t43 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X8 VGND.t80 a_22511_61578# a_22205_61585# VGND.t84 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X9 VGND.t28 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_18252_61704# VGND.t27 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X10 ring_0/inverter_ring_0/skullfet_inverter_6.A ring_0/inverter_ring_0/skullfet_inverter_7.A VDPWR.t29 VDPWR.t28 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X11 VGND.t43 ring_0/inverter_ring_0/skullfet_inverter_13.A ring_0/inverter_ring_0/skullfet_inverter_12.A VGND.t42 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X12 VDPWR.t14 a_20876_61559# a_19955_61640# VDPWR.t2 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X13 a_23109_61717# a_22851_61717# VGND.t13 VGND.t12 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X14 a_24054_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t18 VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X15 VGND.t54 ring_0/inverter_ring_0/skullfet_inverter_17.A ring_0/inverter_ring_0/skullfet_inverter_16.A VGND.t53 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X16 VGND.t26 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_16801_61717# VGND.t25 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X17 a_20876_61559# a_19947_61366# a_20747_61559# VGND.t106 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X18 ring_0/inverter_ring_0/skullfet_inverter_12.A ring_0/inverter_ring_0/skullfet_inverter_13.A VDPWR.t33 VDPWR.t32 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X19 VDPWR.t65 a_22511_61578# freq_divider_0.sg13g2_dfrbp_2_2.D VDPWR.t2 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X20 a_23211_61366# a_23350_61250# VDPWR.t11 VDPWR.t2 sg13_lv_pmos ad=0.3864p pd=2.93u as=1.55707p ps=9.54u w=1.12u l=0.13u
X21 a_23211_61366# a_23350_61250# VGND.t103 VGND.t102 sg13_lv_nmos ad=0.2516p pd=2.16u as=2.07232p ps=13.14u w=0.74u l=0.13u
X22 VGND.t111 ring_0/inverter_ring_0/skullfet_inverter_9.A ring_0/inverter_ring_0/skullfet_inverter_8.A VGND.t110 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X23 ring_0/inverter_ring_0/skullfet_inverter_11.A ring_0/inverter_ring_0/skullfet_inverter_12.A VDPWR.t1 VDPWR.t0 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X24 VDPWR.t34 freq_divider_0.sg13g2_dfrbp_2_2.D a_24054_61326# VDPWR.t2 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X25 a_22851_61717# a_22511_61578# VDPWR.t65 VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X26 a_23161_61402# a_22851_61717# VDPWR.t11 VDPWR.t2 sg13_lv_pmos ad=52.5f pd=0.67u as=1.55707p ps=9.54u w=0.42u l=0.13u
X27 VDPWR.t50 a_16367_61578# a_16061_61585# VDPWR.t2 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X28 a_17996_61559# a_17067_61366# a_17867_61559# VGND.t3 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X29 freq_divider_0.sg13g2_dfrbp_2_1.D a_19247_61578# VDPWR.t68 VDPWR.t2 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X30 VDPWR.t11 a_21777_61520# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t2 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X31 a_22945_61717# a_22511_61578# a_22851_61717# VGND.t83 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X32 VGND.t24 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_24396_61704# VGND.t23 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X33 VDPWR.t63 a_22511_61578# a_22205_61585# VDPWR.t2 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X34 ring_0/inverter_ring_0/skullfet_inverter_3.A ring_0/inverter_ring_0/skullfet_inverter_4.A VDPWR.t8 VDPWR.t7 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X35 a_24396_61704# a_23219_61640# a_24011_61559# VGND.t97 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X36 a_21856_61617# a_21980_61316# VDPWR.t11 VDPWR.t2 sg13_lv_pmos ad=0.2442p pd=2.06u as=1.55707p ps=9.54u w=0.66u l=0.13u
X37 uo_out[2].t1 a_18941_61585# VGND.t61 VGND.t60 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X38 ring_0/inverter_ring_0/skullfet_inverter_17.A ring_0/inverter_ring_0/skullfet_inverter_18.A VDPWR.t60 VDPWR.t59 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X39 VGND.t7 ring_0/inverter_ring_0/skullfet_inverter_14.A ring_0/inverter_ring_0/skullfet_inverter_13.A VGND.t6 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X40 uo_out[2].t0 a_18941_61585# VDPWR.t47 VDPWR.t2 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X41 VGND.t33 ring_0/inverter_ring_0/skullfet_inverter_2.A ring_0/inverter_ring_0/skullfet_inverter_1.A VGND.t32 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X42 a_19247_61578# a_19947_61366# a_19897_61402# VDPWR.t2 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X43 ring_0/inverter_ring_0/skullfet_inverter_4.A ring_0/inverter_ring_0/skullfet_inverter_5.A VDPWR.t25 VDPWR.t24 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X44 VGND.t73 ring_0/inverter_ring_0/skullfet_inverter_11.A ring_0/inverter_ring_0/skullfet_inverter_10.A VGND.t72 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X45 VDPWR.t46 a_18941_61585# uo_out[2].t0 VDPWR.t2 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X46 VGND.t109 ring_0/inverter_ring_0/skullfet_inverter_0.A ring_0/inverter_ring_0/skullfet_inverter_0.Y VGND.t108 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X47 a_20876_61559# a_19947_61366# a_20790_61326# VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X48 a_18106_61326# a_17206_61250# a_17996_61559# VDPWR.t2 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X49 VGND.t41 ring_0/inverter_ring_0/skullfet_inverter_3.A ring_0/inverter_ring_0/skullfet_inverter_2.A VGND.t40 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X50 VGND.t124 ring_0/inverter_ring_0/skullfet_inverter_16.A uo_out[0].t1 VGND.t123 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X51 ring_0/inverter_ring_0/skullfet_inverter_18.A ring_0/inverter_ring_0/skullfet_inverter_19.A VDPWR.t62 VDPWR.t61 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X52 a_19947_61366# a_20086_61250# VDPWR.t11 VDPWR.t2 sg13_lv_pmos ad=0.3864p pd=2.93u as=1.55707p ps=9.54u w=1.12u l=0.13u
X53 ring_0/inverter_ring_0/skullfet_inverter_9.A ring_0/inverter_ring_0/skullfet_inverter_10.A VDPWR.t36 VDPWR.t35 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X54 VGND.t82 a_22511_61578# freq_divider_0.sg13g2_dfrbp_2_2.D VGND.t81 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X55 VGND.t101 uo_out[0].t2 ring_0/inverter_ring_0/skullfet_inverter_14.A VGND.t100 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X56 VGND.t117 a_22205_61585# uo_out[1].t0 VGND.t116 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X57 a_19681_61717# a_19247_61578# a_19587_61717# VGND.t94 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X58 a_17996_61559# a_17067_61366# a_17910_61326# VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X59 a_19955_61640# a_20086_61250# a_19247_61578# VDPWR.t2 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X60 a_20986_61326# a_20086_61250# a_20876_61559# VDPWR.t2 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X61 VDPWR.t12 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_16707_61717# VDPWR.t2 sg13_lv_pmos ad=1.4373p pd=8.805u as=79.8f ps=0.8u w=0.42u l=0.13u
X62 a_24140_61559# a_23211_61366# a_24054_61326# VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X63 a_17067_61366# a_17206_61250# VDPWR.t12 VDPWR.t2 sg13_lv_pmos ad=0.3864p pd=2.93u as=1.55707p ps=9.54u w=1.12u l=0.13u
X64 VDPWR.t11 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_22851_61717# VDPWR.t2 sg13_lv_pmos ad=1.4373p pd=8.805u as=79.8f ps=0.8u w=0.42u l=0.13u
X65 a_17067_61366# a_17206_61250# VGND.t99 VGND.t98 sg13_lv_nmos ad=0.2516p pd=2.16u as=2.07232p ps=13.14u w=0.74u l=0.13u
X66 VDPWR.t45 freq_divider_0.sg13g2_dfrbp_2_0.D a_17910_61326# VDPWR.t2 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X67 freq_divider_0.sg13g2_dfrbp_2_1.D a_19247_61578# VGND.t90 VGND.t93 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X68 a_21132_61704# a_19955_61640# a_20747_61559# VGND.t36 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X69 a_17910_61326# a_17206_61250# a_17996_61559# VGND.t114 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X70 a_19845_61717# a_20086_61250# a_19247_61578# VGND.t88 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X71 a_16965_61717# a_16707_61717# VGND.t26 VGND.t25 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X72 a_19897_61402# a_19587_61717# VDPWR.t12 VDPWR.t2 sg13_lv_pmos ad=52.5f pd=0.67u as=1.55707p ps=9.54u w=0.42u l=0.13u
X73 a_20790_61326# a_20086_61250# a_20876_61559# VGND.t87 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X74 a_18252_61704# a_17075_61640# a_17867_61559# VGND.t74 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X75 VGND.t92 a_19247_61578# freq_divider_0.sg13g2_dfrbp_2_1.D VGND.t91 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X76 VGND.t59 a_18941_61585# uo_out[2].t1 VGND.t58 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X77 a_24140_61559# a_23211_61366# a_24011_61559# VGND.t71 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X78 a_16965_61717# a_17206_61250# a_16367_61578# VGND.t113 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X79 VGND.t90 a_19247_61578# a_18941_61585# VGND.t89 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X80 a_17996_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t13 VDPWR.t2 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X81 VDPWR.t19 a_19955_61640# a_20986_61326# VDPWR.t2 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X82 a_20790_61326# freq_divider_0.sg13g2_dfrbp_2_1.D a_21529_61717# VGND.t52 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X83 VDPWR.t20 a_17996_61559# a_17075_61640# VDPWR.t2 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X84 VGND.t56 ring_0/inverter_ring_0/skullfet_inverter_0.Y ring_0/inverter_ring_0/skullfet_inverter_19.A VGND.t55 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X85 a_24140_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t15 VDPWR.t2 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X86 ring_0/inverter_ring_0/skullfet_inverter_5.A ring_0/inverter_ring_0/skullfet_inverter_6.A VDPWR.t10 VDPWR.t9 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X87 VDPWR.t69 a_19247_61578# freq_divider_0.sg13g2_dfrbp_2_1.D VDPWR.t2 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X88 VGND.t63 ring_0/inverter_ring_0/skullfet_inverter_8.A ring_0/inverter_ring_0/skullfet_inverter_7.A VGND.t62 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X89 VDPWR.t11 uo_out[1].t2 a_20086_61250# VDPWR.t2 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3808p ps=2.92u w=1.12u l=0.13u
X90 VDPWR.t18 a_24140_61559# a_23219_61640# VDPWR.t2 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X91 a_23219_61640# a_23350_61250# a_22511_61578# VDPWR.t2 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X92 VDPWR.t13 a_17075_61640# a_18106_61326# VDPWR.t2 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X93 a_19587_61717# a_19247_61578# VDPWR.t69 VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X94 VGND.t5 ring_0/inverter_ring_0/skullfet_inverter_1.A ring_0/inverter_ring_0/skullfet_inverter_0.A VGND.t4 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X95 ring_0/inverter_ring_0/skullfet_inverter_10.A ring_0/inverter_ring_0/skullfet_inverter_11.A VDPWR.t56 VDPWR.t55 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X96 VDPWR.t86 a_22205_61585# uo_out[1].t1 VDPWR.t2 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X97 VDPWR.t12 uo_out[2].t2 a_17206_61250# VDPWR.t2 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3808p ps=2.92u w=1.12u l=0.13u
X98 VGND.t1 ring_0/inverter_ring_0/skullfet_inverter_12.A ring_0/inverter_ring_0/skullfet_inverter_11.A VGND.t0 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X99 a_23109_61717# a_23350_61250# a_22511_61578# VGND.t121 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X100 ring_0/inverter_ring_0/skullfet_inverter_0.A ring_0/inverter_ring_0/skullfet_inverter_1.A VDPWR.t4 VDPWR.t3 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X101 ring_0/inverter_ring_0/skullfet_inverter_16.A ring_0/inverter_ring_0/skullfet_inverter_17.A VDPWR.t42 VDPWR.t41 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X102 a_21980_61316# a_21980_61316# VGND.t86 VGND.t95 sg13_lv_nmos ad=0.111p pd=1.34u as=2.07232p ps=13.14u w=0.3u l=0.13u
X103 VGND.t22 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_19681_61717# VGND.t21 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X104 ring_0/inverter_ring_0/skullfet_inverter_2.A ring_0/inverter_ring_0/skullfet_inverter_3.A VDPWR.t31 VDPWR.t30 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X105 uo_out[0].t0 ring_0/inverter_ring_0/skullfet_inverter_16.A VDPWR.t89 VDPWR.t88 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X106 a_21529_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t20 VGND.t19 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X107 VGND.t20 a_20876_61559# a_19955_61640# VGND.t31 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X108 uo_out[3].t1 a_16061_61585# VGND.t50 VGND.t49 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X109 VGND.t86 uo_out[1].t2 a_20086_61250# VGND.t85 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.2516p ps=2.16u w=0.74u l=0.13u
X110 VGND.t86 a_21856_61617# a_21777_61520# VGND.t104 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.27427p ps=2.28u w=0.795u l=0.13u
X111 a_16367_61578# a_17067_61366# a_17017_61402# VDPWR.t2 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X112 ring_0/inverter_ring_0/skullfet_inverter_14.A uo_out[0].t2 VDPWR.t77 VDPWR.t76 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X113 VGND.t9 ring_0/inverter_ring_0/skullfet_inverter_4.A ring_0/inverter_ring_0/skullfet_inverter_3.A VGND.t8 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X114 VDPWR.t15 a_23219_61640# a_24250_61326# VDPWR.t2 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X115 a_24250_61326# a_23350_61250# a_24140_61559# VDPWR.t2 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X116 a_20790_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t14 VDPWR.t2 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X117 a_24054_61326# freq_divider_0.sg13g2_dfrbp_2_2.D a_24793_61717# VGND.t44 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X118 a_22511_61578# a_23211_61366# a_23219_61640# VGND.t70 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X119 a_18649_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t18 VGND.t17 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X120 freq_divider_0.sg13g2_dfrbp_2_0.D a_16367_61578# VDPWR.t50 VDPWR.t2 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X121 VGND.t99 uo_out[2].t2 a_17206_61250# VGND.t98 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.2516p ps=2.16u w=0.74u l=0.13u
X122 VDPWR.t68 a_19247_61578# a_18941_61585# VDPWR.t2 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X123 VGND.t39 ring_0/inverter_ring_0/skullfet_inverter_7.A ring_0/inverter_ring_0/skullfet_inverter_6.A VGND.t38 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X124 a_24793_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t16 VGND.t15 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X125 a_17075_61640# a_17206_61250# a_16367_61578# VDPWR.t2 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X126 uo_out[3].t0 a_16061_61585# VDPWR.t38 VDPWR.t2 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X127 a_24054_61326# a_23350_61250# a_24140_61559# VGND.t120 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X128 VDPWR.t37 a_16061_61585# uo_out[3].t0 VDPWR.t2 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X129 a_22511_61578# a_23211_61366# a_23161_61402# VDPWR.t2 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X130 ring_0/inverter_ring_0/skullfet_inverter_8.A ring_0/inverter_ring_0/skullfet_inverter_9.A VDPWR.t82 VDPWR.t81 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X131 uo_out[1].t1 a_22205_61585# VDPWR.t85 VDPWR.t2 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X132 ring_0/inverter_ring_0/skullfet_inverter_7.A ring_0/inverter_ring_0/skullfet_inverter_8.A VDPWR.t49 VDPWR.t48 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X133 VGND.t46 ring_0/inverter_ring_0/skullfet_inverter_10.A ring_0/inverter_ring_0/skullfet_inverter_9.A VGND.t45 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X134 VGND.t16 a_24140_61559# a_23219_61640# VGND.t51 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X135 VGND.t103 uo_out[0].t3 a_23350_61250# VGND.t102 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.2516p ps=2.16u w=0.74u l=0.13u
X136 freq_divider_0.sg13g2_dfrbp_2_2.D a_22511_61578# VDPWR.t63 VDPWR.t2 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X137 a_16801_61717# a_16367_61578# a_16707_61717# VGND.t69 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X138 a_19247_61578# a_19947_61366# a_19955_61640# VGND.t105 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X139 ring_0/inverter_ring_0/skullfet_inverter_1.A ring_0/inverter_ring_0/skullfet_inverter_2.A VDPWR.t23 VDPWR.t22 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X140 ring_0/inverter_ring_0/skullfet_inverter_13.A ring_0/inverter_ring_0/skullfet_inverter_14.A VDPWR.t6 VDPWR.t5 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X141 VDPWR.t12 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_19587_61717# VDPWR.t2 sg13_lv_pmos ad=1.4373p pd=8.805u as=79.8f ps=0.8u w=0.42u l=0.13u
X142 ring_0/inverter_ring_0/skullfet_inverter_0.Y ring_0/inverter_ring_0/skullfet_inverter_0.A VDPWR.t80 VDPWR.t79 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X143 freq_divider_0.sg13g2_dfrbp_2_0.D a_16367_61578# VGND.t65 VGND.t68 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X144 a_17910_61326# freq_divider_0.sg13g2_dfrbp_2_0.D a_18649_61717# VGND.t57 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X145 a_16367_61578# a_17067_61366# a_17075_61640# VGND.t2 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X146 VGND.t13 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_22945_61717# VGND.t12 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X147 a_17017_61402# a_16707_61717# VDPWR.t12 VDPWR.t2 sg13_lv_pmos ad=52.5f pd=0.67u as=1.55707p ps=9.54u w=0.42u l=0.13u
X148 VGND.t76 ring_0/inverter_ring_0/skullfet_inverter_18.A ring_0/inverter_ring_0/skullfet_inverter_17.A VGND.t75 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X149 VGND.t67 a_16367_61578# freq_divider_0.sg13g2_dfrbp_2_0.D VGND.t66 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X150 VGND.t11 ring_0/inverter_ring_0/skullfet_inverter_6.A ring_0/inverter_ring_0/skullfet_inverter_5.A VGND.t10 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X151 VGND.t48 a_16061_61585# uo_out[3].t1 VGND.t47 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X152 a_19845_61717# a_19587_61717# VGND.t22 VGND.t21 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X153 VGND.t35 ring_0/inverter_ring_0/skullfet_inverter_5.A ring_0/inverter_ring_0/skullfet_inverter_4.A VGND.t34 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X154 VGND.t65 a_16367_61578# a_16061_61585# VGND.t64 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X155 VDPWR.t11 uo_out[0].t3 a_23350_61250# VDPWR.t2 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3808p ps=2.92u w=1.12u l=0.13u
X156 a_19947_61366# a_20086_61250# VGND.t86 VGND.t85 sg13_lv_nmos ad=0.2516p pd=2.16u as=2.07232p ps=13.14u w=0.74u l=0.13u
X157 VGND.t78 ring_0/inverter_ring_0/skullfet_inverter_19.A ring_0/inverter_ring_0/skullfet_inverter_18.A VGND.t77 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X158 VDPWR.t40 freq_divider_0.sg13g2_dfrbp_2_1.D a_20790_61326# VDPWR.t2 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X159 freq_divider_0.sg13g2_dfrbp_2_2.D a_22511_61578# VGND.t80 VGND.t79 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
R0 VGND.n202 VGND.n59 36337.9
R1 VGND.n210 VGND.n111 26006.8
R2 VGND.n345 VGND.n111 20289.4
R3 VGND.t8 VGND.n160 19416.2
R4 VGND.n468 VGND.n467 17662.9
R5 VGND.n194 VGND.n70 15262.5
R6 VGND.n202 VGND.n111 12285.4
R7 VGND.n61 VGND.n59 12285.4
R8 VGND.n467 VGND.n466 12279.6
R9 VGND.n200 VGND.t10 12039.2
R10 VGND.t38 VGND.n63 10402.1
R11 VGND.n281 VGND.n274 10052.7
R12 VGND.n469 VGND.n468 10011.4
R13 VGND.n159 VGND.n158 9840.79
R14 VGND.n201 VGND.n61 9066.9
R15 VGND.n265 VGND.n200 7844.55
R16 VGND.n210 VGND.n204 7498.6
R17 VGND.n199 VGND.n198 7474.99
R18 VGND.n158 VGND.n155 7291.79
R19 VGND.n194 VGND.t34 7169.54
R20 VGND.n472 VGND.n65 6899.39
R21 VGND.n476 VGND.n60 6851.13
R22 VGND.n69 VGND.n65 6429.23
R23 VGND.n265 VGND.t40 6051.63
R24 VGND.n203 VGND.n202 6014.02
R25 VGND.n466 VGND.n465 5872.62
R26 VGND.n204 VGND.n203 5699.78
R27 VGND.n466 VGND.n69 5321.16
R28 VGND.n195 VGND.n194 5298.87
R29 VGND.n478 VGND.n477 4953.11
R30 VGND.n468 VGND.n69 4950.06
R31 VGND.n264 VGND.n263 4945.91
R32 VGND.n291 VGND.n155 3511.45
R33 VGND.n158 VGND.n157 3475.34
R34 VGND.n276 VGND.n271 3284.18
R35 VGND.n466 VGND.n71 3154.9
R36 VGND.n200 VGND.n199 3153.12
R37 VGND.n282 VGND.n281 2376.2
R38 VGND.n265 VGND.n157 2220.92
R39 VGND.n470 VGND.n469 2091.57
R40 VGND.n474 VGND.n63 1946.24
R41 VGND.n203 VGND.n201 1880.71
R42 VGND.n160 VGND.n70 1835.32
R43 VGND.n74 VGND.n71 1763.01
R44 VGND.n265 VGND.n201 1734.38
R45 VGND.n200 VGND.n63 1470.05
R46 VGND.n283 VGND.t108 1368.89
R47 VGND.t77 VGND.n276 1347.06
R48 VGND.n276 VGND.t55 1194.61
R49 VGND.t34 VGND.n193 1123.79
R50 VGND.n467 VGND.n70 1061.65
R51 VGND.n283 VGND.n271 977.779
R52 VGND.n60 VGND.t42 964.287
R53 VGND.n265 VGND.n159 905.553
R54 VGND.t42 VGND.n59 876.317
R55 VGND.n476 VGND.n61 837.723
R56 VGND.n275 VGND.n155 814.62
R57 VGND.n237 VGND.n234 744.615
R58 VGND.n486 VGND.n5 744.615
R59 VGND.n53 VGND.n52 744.615
R60 VGND.n209 VGND.t100 675.663
R61 VGND.n198 VGND.t40 656.004
R62 VGND.n465 VGND.t10 656.004
R63 VGND.n199 VGND.t8 615.229
R64 VGND.n159 VGND.n154 608.424
R65 VGND.n346 VGND.n59 575.212
R66 VGND.n199 VGND.n195 498.868
R67 VGND.n237 VGND.t12 480
R68 VGND.n486 VGND.t21 480
R69 VGND.n52 VGND.t25 480
R70 VGND.n471 VGND.t110 455.887
R71 VGND.n74 VGND.t38 427.755
R72 VGND.n265 VGND.n264 402.269
R73 VGND.n477 VGND.n476 395.865
R74 VGND.n265 VGND.n204 392.892
R75 VGND.t6 VGND.n345 372.399
R76 VGND.n282 VGND.n271 344.149
R77 VGND.t55 VGND.n274 335.173
R78 VGND.n68 VGND.t110 330.428
R79 VGND.n291 VGND.t53 318.406
R80 VGND.n345 VGND.n344 307.757
R81 VGND.n160 VGND.n157 278.079
R82 VGND.n233 VGND.t81 260.005
R83 VGND.n16 VGND.t91 260.005
R84 VGND.t66 VGND.n54 260.005
R85 VGND.t79 VGND.n231 234.738
R86 VGND.t93 VGND.n14 234.738
R87 VGND.n56 VGND.t68 234.738
R88 VGND.n244 VGND.t84 232.869
R89 VGND.n25 VGND.t89 232.869
R90 VGND.t64 VGND.n43 232.869
R91 VGND.t32 VGND.n154 231.615
R92 VGND.t104 VGND.n228 228.233
R93 VGND.n275 VGND.t4 227.947
R94 VGND.n201 VGND.n63 226.054
R95 VGND.n251 VGND.t31 200.339
R96 VGND.n31 VGND.t37 200.339
R97 VGND.n215 VGND.t51 200.339
R98 VGND.n249 VGND.t52 195.942
R99 VGND.n12 VGND.t57 194.969
R100 VGND.n475 VGND.n474 194.851
R101 VGND.n248 VGND.t116 185.124
R102 VGND.n29 VGND.t58 185.124
R103 VGND.t47 VGND.n41 185.124
R104 VGND.t118 VGND.n229 184.825
R105 VGND.t60 VGND.n12 184.825
R106 VGND.n263 VGND.t44 180.052
R107 VGND.n229 VGND.t95 172.145
R108 VGND.n478 VGND.t49 169.907
R109 VGND.n281 VGND.t75 164.255
R110 VGND.t36 VGND.t29 159.763
R111 VGND.t74 VGND.t27 159.763
R112 VGND.t97 VGND.t23 159.763
R113 VGND.t106 VGND.n224 156.929
R114 VGND.t3 VGND.n9 156.929
R115 VGND.t71 VGND.n212 156.929
R116 VGND.n255 VGND.t87 154.614
R117 VGND.n35 VGND.t114 154.614
R118 VGND.n218 VGND.t120 154.614
R119 VGND.n71 VGND.n65 151.276
R120 VGND.t19 VGND.n226 149.62
R121 VGND.t17 VGND.n11 149.62
R122 VGND.t15 VGND.n214 149.62
R123 VGND.t12 VGND.t70 138.463
R124 VGND.t21 VGND.t105 138.463
R125 VGND.t25 VGND.t2 138.463
R126 VGND.n264 VGND.t123 132.323
R127 VGND.n474 VGND.t62 128.216
R128 VGND.n477 VGND.n59 122.921
R129 VGND.t108 VGND.n282 113.026
R130 VGND.n234 VGND.t83 110.237
R131 VGND.t94 VGND.n5 110.237
R132 VGND.t69 VGND.n53 110.237
R133 VGND.n224 VGND.n5 106.212
R134 VGND.n53 VGND.n9 106.212
R135 VGND.n234 VGND.n212 106.212
R136 VGND.t87 VGND.n254 100.478
R137 VGND.t114 VGND.n34 100.478
R138 VGND.t120 VGND.n217 100.478
R139 VGND.n255 VGND.t106 99.7516
R140 VGND.n35 VGND.t3 99.7516
R141 VGND.n218 VGND.t71 99.7516
R142 VGND.n469 VGND.n68 95.8456
R143 VGND.t62 VGND.n473 95.5275
R144 VGND.n251 VGND.t19 93.8297
R145 VGND.n31 VGND.t17 93.8297
R146 VGND.n215 VGND.t15 93.8297
R147 VGND.t95 VGND.n228 86.222
R148 VGND.n291 VGND.n154 84.6642
R149 VGND.n473 VGND.n472 83.8532
R150 VGND.n254 VGND.t36 75.5501
R151 VGND.n34 VGND.t74 75.5501
R152 VGND.n217 VGND.t97 75.5501
R153 VGND.t102 VGND.t121 73.8467
R154 VGND.t85 VGND.t88 73.8467
R155 VGND.t98 VGND.t113 73.8467
R156 VGND.n248 VGND.t118 73.5423
R157 VGND.n29 VGND.t60 73.5423
R158 VGND.t49 VGND.n41 73.5423
R159 VGND.t116 VGND.n244 73.244
R160 VGND.t58 VGND.n25 73.244
R161 VGND.n43 VGND.t47 73.244
R162 VGND.n290 VGND.t4 72.396
R163 VGND.n344 VGND.t100 65.0575
R164 VGND.n346 VGND.t6 63.8663
R165 VGND.n476 VGND.t0 63.5677
R166 VGND.t52 VGND.n226 63.3986
R167 VGND.t57 VGND.n11 63.3986
R168 VGND.n214 VGND.t44 63.3986
R169 VGND.t51 VGND.n213 59.0031
R170 VGND.t31 VGND.n225 59.0031
R171 VGND.t37 VGND.n10 59.0031
R172 VGND.n474 VGND.t72 55.0827
R173 VGND.n266 VGND.t32 51.425
R174 VGND.n206 VGND.t53 51.1311
R175 VGND.t83 VGND.n233 48.4827
R176 VGND.n16 VGND.t94 48.4827
R177 VGND.n54 VGND.t69 48.4827
R178 VGND.t0 VGND.n475 47.9255
R179 VGND.n471 VGND.t45 47.7166
R180 VGND.n471 VGND.n66 44.7738
R181 VGND.n292 VGND.t75 44.7032
R182 VGND.t123 VGND.n210 42.4247
R183 VGND.n66 VGND.t72 41.6077
R184 VGND.n280 VGND.t77 38.7252
R185 VGND.t29 VGND.n225 38.7147
R186 VGND.t27 VGND.n10 38.7147
R187 VGND.t23 VGND.n213 38.7147
R188 VGND.n281 VGND.n275 36.6123
R189 VGND.t45 VGND.n470 36.1063
R190 VGND.n249 VGND.t104 31.1079
R191 VGND.t84 VGND.n231 28.3754
R192 VGND.t89 VGND.n14 28.3754
R193 VGND.n56 VGND.t64 28.3754
R194 VGND.n232 VGND.t79 27.8464
R195 VGND.n15 VGND.t93 27.8464
R196 VGND.t68 VGND.n55 27.8464
R197 VGND.t70 VGND.t102 24.6159
R198 VGND.t105 VGND.t85 24.6159
R199 VGND.t2 VGND.t98 24.6159
R200 VGND.n291 VGND.n290 22.6588
R201 VGND.n210 VGND.n209 22.6333
R202 VGND.n472 VGND.n471 18.8055
R203 VGND.n289 VGND.n288 18.1658
R204 VGND.n268 VGND.n267 18.1658
R205 VGND.n88 VGND.n62 18.1658
R206 VGND.n393 VGND.n392 18.1658
R207 VGND.n77 VGND.n64 18.1658
R208 VGND.n76 VGND.n75 18.1658
R209 VGND.n464 VGND.n463 18.1658
R210 VGND.n193 VGND.n192 18.1658
R211 VGND.n162 VGND.n161 18.1658
R212 VGND.n448 VGND.n447 18.1658
R213 VGND.n87 VGND.n67 18.1658
R214 VGND.n208 VGND.n207 18.1658
R215 VGND.n294 VGND.n293 18.1658
R216 VGND.n279 VGND.n278 18.1658
R217 VGND.n273 VGND.n272 18.1658
R218 VGND.n205 VGND.n141 18.1658
R219 VGND.n343 VGND.n342 18.1658
R220 VGND.n348 VGND.n347 18.1658
R221 VGND.n374 VGND.n373 18.1658
R222 VGND.n197 VGND.n196 18.1658
R223 VGND.n285 VGND.n284 18.1658
R224 VGND.t86 VGND.n255 18.0261
R225 VGND.t99 VGND.n35 18.0261
R226 VGND.t103 VGND.n218 18.0261
R227 VGND.t81 VGND.n232 17.5282
R228 VGND.t91 VGND.n15 17.5282
R229 VGND.n55 VGND.t66 17.5282
R230 VGND.n216 VGND.t16 17.2928
R231 VGND.n36 VGND.t28 17.2395
R232 VGND.n256 VGND.t30 17.2395
R233 VGND.n219 VGND.t24 17.2395
R234 VGND.n47 VGND.t67 17.2297
R235 VGND.n21 VGND.t92 17.2297
R236 VGND.n240 VGND.t82 17.2297
R237 VGND.n40 VGND.t26 17.2268
R238 VGND.n32 VGND.t18 17.2268
R239 VGND.n19 VGND.t22 17.2268
R240 VGND.n252 VGND.t20 17.2268
R241 VGND.n223 VGND.t13 17.2268
R242 VGND.n404 VGND.t65 17.212
R243 VGND.n23 VGND.t90 17.212
R244 VGND.n242 VGND.t80 17.212
R245 VGND.n57 VGND.t50 17.2025
R246 VGND.n27 VGND.t61 17.2025
R247 VGND.n246 VGND.t119 17.2025
R248 VGND.n289 VGND.t5 17.0362
R249 VGND.n267 VGND.t33 17.0362
R250 VGND.n62 VGND.t1 17.0362
R251 VGND.n392 VGND.t73 17.0362
R252 VGND.n64 VGND.t63 17.0362
R253 VGND.n75 VGND.t39 17.0362
R254 VGND.n464 VGND.t11 17.0362
R255 VGND.n193 VGND.t35 17.0362
R256 VGND.n161 VGND.t9 17.0362
R257 VGND.n447 VGND.t111 17.0362
R258 VGND.n67 VGND.t46 17.0362
R259 VGND.n208 VGND.t124 17.0362
R260 VGND.n293 VGND.t76 17.0362
R261 VGND.n279 VGND.t78 17.0362
R262 VGND.n273 VGND.t56 17.0362
R263 VGND.n205 VGND.t54 17.0362
R264 VGND.n343 VGND.t101 17.0362
R265 VGND.n347 VGND.t7 17.0362
R266 VGND.n373 VGND.t43 17.0362
R267 VGND.n197 VGND.t41 17.0362
R268 VGND.n284 VGND.t109 17.0362
R269 VGND.n263 VGND.t103 17.0005
R270 VGND.t103 VGND.n214 17.0005
R271 VGND.t103 VGND.n215 17.0005
R272 VGND.n258 VGND.t86 17.0005
R273 VGND.t86 VGND.n231 17.0005
R274 VGND.t86 VGND.n248 17.0005
R275 VGND.t86 VGND.n230 17.0005
R276 VGND.t86 VGND.n228 17.0005
R277 VGND.t86 VGND.n226 17.0005
R278 VGND.t86 VGND.n251 17.0005
R279 VGND.n488 VGND.n1 17.0005
R280 VGND.n489 VGND.n488 17.0005
R281 VGND.t99 VGND.n18 17.0005
R282 VGND.t99 VGND.n14 17.0005
R283 VGND.t99 VGND.n29 17.0005
R284 VGND.t99 VGND.n13 17.0005
R285 VGND.t99 VGND.n11 17.0005
R286 VGND.t99 VGND.n31 17.0005
R287 VGND.n480 VGND.n479 17.0005
R288 VGND.n479 VGND.n56 17.0005
R289 VGND.n479 VGND.n41 17.0005
R290 VGND.n479 VGND.n58 17.0005
R291 VGND.n479 VGND.n478 17.0005
R292 VGND.n284 VGND.n283 16.9935
R293 VGND.n266 VGND.n265 16.2915
R294 VGND.n265 VGND.n206 16.2014
R295 VGND.n470 VGND.n67 15.6652
R296 VGND.n280 VGND.n279 15.5838
R297 VGND.n392 VGND.n66 15.4962
R298 VGND.n293 VGND.n292 15.4044
R299 VGND.n475 VGND.n62 15.3111
R300 VGND.n206 VGND.n205 15.2207
R301 VGND.n267 VGND.n266 15.2126
R302 VGND.n347 VGND.n346 14.8829
R303 VGND.n209 VGND.n208 14.853
R304 VGND.n344 VGND.n343 14.853
R305 VGND.n290 VGND.n289 14.6742
R306 VGND.n292 VGND.n291 14.2225
R307 VGND.n473 VGND.n64 14.1685
R308 VGND.n281 VGND.n280 12.3693
R309 VGND.n491 VGND.n490 11.5981
R310 VGND.n406 VGND.n405 11.5903
R311 VGND.n447 VGND.n68 11.5621
R312 VGND.n274 VGND.n273 11.5336
R313 VGND.n75 VGND.n74 11.0666
R314 VGND.n465 VGND.n464 10.3577
R315 VGND.n198 VGND.n197 10.3577
R316 VGND.n373 VGND.n60 9.85117
R317 VGND.n195 VGND.n161 9.69267
R318 VGND.n435 VGND.n430 9.0005
R319 VGND.n430 VGND.n423 9.0005
R320 VGND.n435 VGND.n434 9.0005
R321 VGND.n434 VGND.n423 9.0005
R322 VGND.n435 VGND.n429 9.0005
R323 VGND.n436 VGND.n425 9.0005
R324 VGND.n436 VGND.n423 9.0005
R325 VGND.n436 VGND.n435 9.0005
R326 VGND.n441 VGND.n438 9.0005
R327 VGND.n438 VGND.n421 9.0005
R328 VGND.n441 VGND.n440 9.0005
R329 VGND.n440 VGND.n421 9.0005
R330 VGND.n441 VGND.n437 9.0005
R331 VGND.n443 VGND.n442 9.0005
R332 VGND.n442 VGND.n421 9.0005
R333 VGND.n442 VGND.n441 9.0005
R334 VGND.n442 uio_oe[7] 8.8478
R335 VGND.n44 VGND.t48 8.74885
R336 VGND.n26 VGND.t59 8.74885
R337 VGND.n245 VGND.t117 8.74885
R338 VGND.n237 VGND.n235 8.501
R339 VGND.n237 VGND.n236 8.501
R340 VGND.n487 VGND.n486 8.501
R341 VGND.n486 VGND.n6 8.501
R342 VGND.n52 VGND.n50 8.501
R343 VGND.n52 VGND.n51 8.501
R344 VGND.n261 VGND.n220 8.47111
R345 VGND.n260 VGND.n221 8.47111
R346 VGND.n259 VGND.n222 8.47111
R347 VGND.t86 VGND.n241 8.47111
R348 VGND.t86 VGND.n243 8.47111
R349 VGND.t86 VGND.n247 8.47111
R350 VGND.t86 VGND.n253 8.47111
R351 VGND.n4 VGND.n2 8.47111
R352 VGND.n17 VGND.n7 8.47111
R353 VGND.t99 VGND.n22 8.47111
R354 VGND.t99 VGND.n24 8.47111
R355 VGND.t99 VGND.n28 8.47111
R356 VGND.t99 VGND.n33 8.47111
R357 VGND.n483 VGND.n37 8.47111
R358 VGND.n482 VGND.n38 8.47111
R359 VGND.n481 VGND.n39 8.47111
R360 VGND.n479 VGND.n46 8.47111
R361 VGND.n479 VGND.n45 8.47111
R362 VGND.n479 VGND.n42 8.47111
R363 VGND.n269 VGND.n156 8.0799
R364 VGND.n460 VGND.n459 7.52168
R365 VGND.n460 VGND.n76 7.47272
R366 VGND.n277 VGND.n153 6.68645
R367 VGND.n394 VGND.n391 6.63864
R368 VGND.n463 VGND.n462 6.53659
R369 VGND.n163 VGND.n162 6.32858
R370 VGND.n192 VGND.n191 6.07977
R371 VGND.n196 VGND.n156 6.05718
R372 VGND.n269 VGND.n268 5.9638
R373 VGND.n238 VGND.n237 5.66778
R374 VGND.n486 VGND.n485 5.66778
R375 VGND.n52 VGND.n49 5.66778
R376 VGND.n237 VGND.n211 5.66767
R377 VGND.n486 VGND.n3 5.66767
R378 VGND.n52 VGND.n8 5.66767
R379 VGND.t86 VGND.n239 5.61485
R380 VGND.t86 VGND.n250 5.61485
R381 VGND.t99 VGND.n20 5.61485
R382 VGND.t99 VGND.n30 5.61485
R383 VGND.n479 VGND.n48 5.61485
R384 VGND.n287 VGND.n269 5.51412
R385 VGND.n429 VGND 5.4103
R386 VGND.n288 VGND.n287 4.6955
R387 VGND.n433 VGND.n432 4.49573
R388 VGND.n432 VGND.n424 4.49573
R389 VGND.n439 VGND.n396 4.49573
R390 VGND.n422 VGND.n396 4.49573
R391 VGND.n431 VGND.n425 4.49573
R392 VGND.n443 VGND.n399 4.49573
R393 VGND.n429 VGND.n428 4.4949
R394 VGND.n437 VGND.n398 4.4949
R395 VGND.n286 VGND.n285 4.09378
R396 VGND.n272 VGND.n270 3.42765
R397 VGND.t103 VGND.n216 3.38768
R398 VGND.t86 VGND.n227 3.34182
R399 VGND.n278 VGND.n277 3.27628
R400 VGND.n295 VGND.n294 2.85446
R401 VGND.n322 VGND.n125 2.31911
R402 VGND.n125 VGND 2.31911
R403 VGND.n78 VGND.n77 2.27849
R404 VGND.n445 VGND.n396 2.2505
R405 VGND.n444 VGND.n443 2.2505
R406 VGND.n432 VGND.n86 2.2505
R407 VGND.n426 VGND.n425 2.2505
R408 VGND.t103 VGND.n262 1.97699
R409 VGND.t86 VGND.n257 1.97699
R410 VGND.t99 VGND.n484 1.97699
R411 VGND.n307 VGND.n141 1.86972
R412 VGND.n449 VGND.n448 1.81263
R413 VGND.n342 VGND.n341 1.47805
R414 VGND.n341 VGND.n340 1.4745
R415 VGND.n395 VGND.n87 1.41597
R416 VGND.n437 VGND.n436 1.40696
R417 VGND.t86 VGND.n254 1.21402
R418 VGND.t99 VGND.n34 1.21402
R419 VGND.t103 VGND.n217 1.21402
R420 VGND.n277 VGND.n270 1.18201
R421 VGND.n444 VGND.n397 1.1463
R422 VGND.n427 VGND.n426 1.1463
R423 VGND.n394 VGND.n393 1.13055
R424 VGND.n89 VGND.n88 1.1093
R425 VGND.t103 VGND.n212 1.04263
R426 VGND.t86 VGND.n244 1.04263
R427 VGND.t86 VGND.n229 1.04263
R428 VGND.t86 VGND.n224 1.04263
R429 VGND.t99 VGND.n25 1.04263
R430 VGND.t99 VGND.n12 1.04263
R431 VGND.t99 VGND.n9 1.04263
R432 VGND.n479 VGND.n43 1.04263
R433 VGND.t86 VGND.n233 1.02715
R434 VGND.t86 VGND.n232 1.02715
R435 VGND.t99 VGND.n16 1.02715
R436 VGND.t99 VGND.n15 1.02715
R437 VGND.n479 VGND.n54 1.02715
R438 VGND.n479 VGND.n55 1.02715
R439 VGND.n324 VGND.n125 0.936079
R440 VGND.n207 VGND.n125 0.851167
R441 VGND.n349 VGND.n348 0.8068
R442 VGND.n375 VGND.n374 0.803036
R443 VGND.n395 VGND.n394 0.610292
R444 VGND.n379 VGND.n378 0.598489
R445 VGND.n307 VGND.n306 0.597922
R446 VGND.n262 VGND.n261 0.585769
R447 VGND.n484 VGND.n483 0.585769
R448 VGND.n257 VGND.n1 0.52548
R449 VGND.n446 VGND.n445 0.521717
R450 VGND.n461 VGND.n460 0.518224
R451 VGND.n262 VGND.n219 0.477006
R452 VGND.n257 VGND.n256 0.477006
R453 VGND.n484 VGND.n36 0.477006
R454 VGND.n341 VGND.n112 0.473781
R455 VGND.n163 VGND.n156 0.464095
R456 VGND.n451 VGND.n86 0.45348
R457 VGND.n337 VGND.n112 0.434656
R458 VGND.n380 VGND.n379 0.352948
R459 VGND.n306 VGND.n305 0.352948
R460 VGND.n337 VGND.n336 0.347746
R461 VGND.n164 VGND.n163 0.328048
R462 VGND.n287 VGND.n286 0.326045
R463 VGND.n400 uo_out[5] 0.32522
R464 VGND.n401 uo_out[6] 0.32522
R465 VGND.n402 uo_out[7] 0.32522
R466 VGND.n403 uio_out[0] 0.32522
R467 VGND.n408 uio_out[2] 0.32522
R468 VGND.n409 uio_out[3] 0.32522
R469 VGND.n410 uio_out[4] 0.32522
R470 VGND.n411 uio_out[5] 0.32522
R471 VGND.n412 uio_out[6] 0.32522
R472 VGND.n413 uio_out[7] 0.32522
R473 VGND.n414 uio_oe[0] 0.32522
R474 VGND.n415 uio_oe[1] 0.32522
R475 VGND.n416 uio_oe[2] 0.32522
R476 VGND.n417 uio_oe[3] 0.32522
R477 VGND.n418 uio_oe[4] 0.32522
R478 VGND.n419 uio_oe[5] 0.32522
R479 VGND.n420 uio_oe[6] 0.32522
R480 VGND.n336 VGND.n335 0.289181
R481 VGND.n491 VGND.n0 0.27022
R482 VGND.n381 VGND.n380 0.2683
R483 VGND.n305 VGND.n304 0.2683
R484 VGND.n189 VGND.n164 0.256021
R485 VGND.n340 VGND.n110 0.250193
R486 VGND.n449 VGND.n446 0.243514
R487 VGND.n335 VGND.n334 0.243383
R488 VGND VGND.n227 0.243171
R489 VGND.n261 VGND.n260 0.241078
R490 VGND.n260 VGND.n259 0.241078
R491 VGND.n17 VGND.n2 0.241078
R492 VGND.n483 VGND.n482 0.241078
R493 VGND.n482 VGND.n481 0.241078
R494 VGND VGND.n227 0.237591
R495 VGND.n407 VGND.n406 0.22226
R496 VGND.n382 VGND.n381 0.221084
R497 VGND.n304 VGND.n303 0.221084
R498 VGND.n334 VGND.n333 0.216589
R499 VGND.n219 VGND.n216 0.208
R500 VGND.n286 VGND.n270 0.201227
R501 VGND.n383 VGND.n382 0.193014
R502 VGND.n303 VGND.n302 0.193014
R503 VGND.n333 VGND.n332 0.189923
R504 VGND.n250 VGND 0.180825
R505 VGND.n30 VGND 0.180825
R506 VGND.n259 VGND.n258 0.180789
R507 VGND.n489 VGND.n2 0.180789
R508 VGND.n18 VGND.n17 0.180789
R509 VGND.n481 VGND.n480 0.180789
R510 VGND.n240 VGND.n239 0.177986
R511 VGND.n21 VGND.n20 0.177986
R512 VGND.n48 VGND.n47 0.177986
R513 VGND.n332 VGND.n331 0.177878
R514 VGND.n384 VGND.n383 0.172356
R515 VGND.n302 VGND.n301 0.172356
R516 VGND.n189 VGND.n188 0.165165
R517 VGND.n253 VGND.n252 0.163289
R518 VGND.n33 VGND.n32 0.163289
R519 VGND.n331 VGND.n330 0.161737
R520 VGND.n247 VGND.n246 0.159539
R521 VGND.n28 VGND.n27 0.159539
R522 VGND.n57 VGND.n42 0.159539
R523 VGND.n461 VGND.n73 0.158526
R524 VGND.n239 VGND.n223 0.158325
R525 VGND.n20 VGND.n19 0.158325
R526 VGND.n48 VGND.n40 0.158325
R527 VGND.n385 VGND.n384 0.155671
R528 VGND.n301 VGND.n300 0.155671
R529 VGND.n188 VGND.n187 0.152148
R530 VGND.n390 VGND.n389 0.150927
R531 VGND.n330 VGND.n329 0.149148
R532 VGND.n388 VGND.n90 0.149023
R533 VGND.n387 VGND.n91 0.147167
R534 VGND.n298 VGND.n150 0.147167
R535 VGND.n187 VGND.n186 0.145833
R536 VGND.n245 VGND.n243 0.145789
R537 VGND.n26 VGND.n24 0.145789
R538 VGND.n45 VGND.n44 0.145789
R539 VGND.n386 VGND.n92 0.144762
R540 VGND.n299 VGND.n149 0.144762
R541 VGND.n386 VGND.n385 0.143511
R542 VGND.n300 VGND.n299 0.143511
R543 VGND.n153 VGND.n152 0.143335
R544 VGND.n385 VGND.n93 0.14301
R545 VGND.n300 VGND.n148 0.14301
R546 VGND.n329 VGND.n328 0.142866
R547 VGND.n384 VGND.n94 0.1413
R548 VGND.n301 VGND.n147 0.1413
R549 VGND.n383 VGND.n95 0.13963
R550 VGND.n302 VGND.n146 0.13963
R551 VGND.n391 VGND.n89 0.139117
R552 VGND.n382 VGND.n96 0.138
R553 VGND.n303 VGND.n145 0.138
R554 VGND.n252 VGND.n250 0.137986
R555 VGND.n32 VGND.n30 0.137986
R556 VGND.n186 VGND.n185 0.136464
R557 VGND.n381 VGND.n97 0.136407
R558 VGND.n304 VGND.n144 0.136407
R559 VGND.n456 VGND.n455 0.134991
R560 VGND.n380 VGND.n98 0.134851
R561 VGND.n305 VGND.n143 0.134851
R562 VGND.n387 VGND.n386 0.134721
R563 VGND.n299 VGND.n298 0.134721
R564 VGND.n328 VGND.n327 0.133592
R565 VGND.n379 VGND.n99 0.13333
R566 VGND.n306 VGND.n142 0.13333
R567 VGND.n185 VGND.n184 0.131588
R568 VGND.n242 VGND.n241 0.130789
R569 VGND.n23 VGND.n22 0.130789
R570 VGND.n327 VGND.n326 0.127631
R571 VGND.n350 VGND.n109 0.127631
R572 VGND.n388 VGND.n387 0.127467
R573 VGND.n298 VGND.n297 0.127467
R574 VGND.n184 VGND.n183 0.126098
R575 VGND.n326 VGND.n325 0.123294
R576 VGND.n241 VGND.n240 0.123289
R577 VGND.n22 VGND.n21 0.123289
R578 VGND.n47 VGND.n46 0.123289
R579 VGND.n354 VGND.n109 0.122221
R580 VGND.n349 VGND.n110 0.122211
R581 VGND.n183 VGND.n182 0.121629
R582 VGND.n389 VGND.n388 0.121573
R583 VGND.n297 VGND.n296 0.121573
R584 VGND.n405 VGND.n46 0.120789
R585 VGND.n391 VGND.n390 0.119995
R586 VGND.n177 VGND.n176 0.119457
R587 VGND.n182 VGND.n181 0.118673
R588 VGND.n355 VGND.n354 0.117844
R589 VGND.n177 VGND.n73 0.117211
R590 VGND.n181 VGND.n180 0.114913
R591 VGND.n356 VGND.n355 0.114675
R592 VGND.n180 VGND.n179 0.113743
R593 VGND.n339 VGND.n112 0.112734
R594 VGND.n338 VGND.n337 0.112578
R595 VGND.n256 VGND.n253 0.112039
R596 VGND.n36 VGND.n33 0.112039
R597 VGND.n336 VGND.n113 0.111718
R598 VGND.n335 VGND.n114 0.111507
R599 VGND.n321 VGND.n320 0.111202
R600 VGND.n356 VGND.n107 0.111202
R601 VGND.n297 VGND.n151 0.11115
R602 VGND.n243 VGND.n242 0.110789
R603 VGND.n24 VGND.n23 0.110789
R604 VGND.n404 VGND.n45 0.110789
R605 VGND.n179 VGND.n178 0.110741
R606 VGND.n334 VGND.n115 0.110644
R607 VGND.n178 VGND.n177 0.110231
R608 VGND.n333 VGND.n116 0.110139
R609 VGND.n320 VGND.n319 0.110119
R610 VGND.n332 VGND.n117 0.109632
R611 VGND.n190 VGND.n189 0.109257
R612 VGND.n360 VGND.n107 0.109256
R613 VGND.n331 VGND.n118 0.109053
R614 VGND.n188 VGND.n165 0.10874
R615 VGND.n330 VGND.n119 0.10854
R616 VGND.n187 VGND.n166 0.108513
R617 VGND.n186 VGND.n167 0.108352
R618 VGND.n185 VGND.n168 0.108122
R619 VGND.n329 VGND.n120 0.108023
R620 VGND.n328 VGND.n121 0.107796
R621 VGND.n183 VGND.n170 0.107722
R622 VGND.n184 VGND.n169 0.107592
R623 VGND.n182 VGND.n171 0.107552
R624 VGND.n180 VGND.n173 0.10751
R625 VGND.n327 VGND.n122 0.107273
R626 VGND.n351 VGND.n350 0.107273
R627 VGND.n319 VGND.n318 0.107182
R628 VGND.n178 VGND.n175 0.107092
R629 VGND.n326 VGND.n123 0.107042
R630 VGND.n352 VGND.n109 0.107042
R631 VGND.n181 VGND.n172 0.10701
R632 VGND.n179 VGND.n174 0.106962
R633 VGND.n325 VGND.n124 0.10687
R634 VGND.n354 VGND.n353 0.10687
R635 VGND.n323 VGND.n126 0.106635
R636 VGND.n355 VGND.n108 0.106635
R637 VGND.n377 VGND.n101 0.106426
R638 VGND.n309 VGND.n139 0.106426
R639 VGND.n361 VGND.n360 0.106367
R640 VGND.n321 VGND.n127 0.1061
R641 VGND.n357 VGND.n356 0.1061
R642 VGND.n319 VGND.n129 0.10604
R643 VGND.n360 VGND.n359 0.10604
R644 VGND.n317 VGND.n131 0.105977
R645 VGND.n363 VGND.n362 0.105977
R646 VGND.n312 VGND.n136 0.105973
R647 VGND.n370 VGND.n103 0.105973
R648 VGND.n320 VGND.n128 0.10592
R649 VGND.n358 VGND.n107 0.10592
R650 VGND.n376 VGND.n102 0.105907
R651 VGND.n310 VGND.n138 0.105907
R652 VGND.n313 VGND.n135 0.105848
R653 VGND.n369 VGND.n368 0.105848
R654 VGND.n311 VGND.n137 0.10578
R655 VGND.n372 VGND.n371 0.10578
R656 VGND.n316 VGND.n132 0.105731
R657 VGND.n364 VGND.n105 0.105731
R658 VGND.n318 VGND.n317 0.105665
R659 VGND.n314 VGND.n134 0.105663
R660 VGND.n367 VGND.n104 0.105663
R661 VGND.n315 VGND.n133 0.105542
R662 VGND.n366 VGND.n365 0.105542
R663 VGND.n318 VGND.n130 0.105493
R664 VGND.n361 VGND.n106 0.105493
R665 VGND.n362 VGND.n361 0.104886
R666 VGND.n295 VGND.n153 0.104495
R667 VGND.n317 VGND.n316 0.104166
R668 VGND.n362 VGND.n105 0.104166
R669 VGND.n406 uio_out[1] 0.10346
R670 VGND.n315 VGND.n314 0.102551
R671 VGND.n316 VGND.n315 0.102053
R672 VGND.n366 VGND.n105 0.102053
R673 VGND.n322 VGND.n321 0.101891
R674 VGND.n367 VGND.n366 0.101858
R675 VGND.n314 VGND.n313 0.101493
R676 VGND.n368 VGND.n367 0.101493
R677 VGND.n313 VGND.n312 0.100967
R678 VGND.n368 VGND.n103 0.100967
R679 VGND.n310 VGND.n309 0.100958
R680 VGND.n311 VGND.n310 0.100445
R681 VGND.n377 VGND.n376 0.100376
R682 VGND.n312 VGND.n311 0.100187
R683 VGND.n372 VGND.n103 0.100187
R684 VGND.n73 VGND.n72 0.0973571
R685 VGND.n247 VGND.n245 0.095789
R686 VGND.n28 VGND.n26 0.095789
R687 VGND.n44 VGND.n42 0.095789
R688 VGND.n455 VGND.n454 0.0954338
R689 VGND.n450 VGND.n85 0.0928432
R690 VGND.n325 VGND.n324 0.0895217
R691 VGND.n459 VGND.n458 0.0873393
R692 VGND.n207 VGND 0.0854123
R693 VGND.n258 VGND.n223 0.083
R694 VGND.n19 VGND.n18 0.083
R695 VGND.n480 VGND.n40 0.083
R696 VGND.n378 VGND.n100 0.0802603
R697 VGND.n308 VGND.n140 0.0802603
R698 VGND.n101 VGND.n100 0.0782828
R699 VGND.n140 VGND.n139 0.0782828
R700 VGND.n490 VGND.n489 0.078
R701 VGND.n390 VGND.n90 0.0779701
R702 VGND.n376 VGND.n375 0.0771258
R703 VGND.n350 VGND.n349 0.0762778
R704 VGND.n454 VGND.n453 0.0754235
R705 VGND.n91 VGND.n90 0.0751329
R706 VGND.n450 VGND.n449 0.0739655
R707 VGND.n151 VGND.n150 0.0735315
R708 VGND.n92 VGND.n91 0.0731
R709 VGND.n150 VGND.n149 0.0731
R710 VGND.n458 VGND.n79 0.0724725
R711 VGND.n93 VGND.n92 0.0701066
R712 VGND.n149 VGND.n148 0.0701066
R713 VGND.n94 VGND.n93 0.067836
R714 VGND.n148 VGND.n147 0.067836
R715 VGND.n95 VGND.n94 0.06562
R716 VGND.n147 VGND.n146 0.06562
R717 VGND.t103 VGND.n213 0.0650946
R718 VGND.t86 VGND.n249 0.0650946
R719 VGND.t86 VGND.n225 0.0650946
R720 VGND.t99 VGND.n10 0.0650946
R721 VGND.n96 VGND.n95 0.0634565
R722 VGND.n146 VGND.n145 0.0634565
R723 VGND.n453 VGND.n452 0.0614573
R724 VGND.n288 VGND 0.061
R725 VGND.n268 VGND 0.061
R726 VGND.n393 VGND 0.061
R727 VGND.n77 VGND 0.061
R728 VGND.n76 VGND 0.061
R729 VGND.n463 VGND 0.061
R730 VGND.n192 VGND 0.061
R731 VGND.n162 VGND 0.061
R732 VGND.n448 VGND 0.061
R733 VGND.n87 VGND 0.061
R734 VGND.n88 VGND 0.061
R735 VGND.n97 VGND.n96 0.061
R736 VGND.n294 VGND 0.061
R737 VGND.n278 VGND 0.061
R738 VGND.n272 VGND 0.061
R739 VGND.n145 VGND.n144 0.061
R740 VGND.n141 VGND 0.061
R741 VGND.n342 VGND 0.061
R742 VGND.n348 VGND 0.061
R743 VGND.n374 VGND 0.061
R744 VGND.n196 VGND 0.061
R745 VGND.n285 VGND 0.061
R746 VGND.n81 VGND.n80 0.0607651
R747 VGND.n230 VGND 0.0605
R748 VGND VGND.n13 0.0605
R749 VGND.n58 VGND 0.0605
R750 VGND.n98 VGND.n97 0.0589402
R751 VGND.n144 VGND.n143 0.0589402
R752 VGND.n452 VGND.n451 0.0585315
R753 VGND.n296 VGND.n152 0.0568276
R754 VGND.n99 VGND.n98 0.0565916
R755 VGND.n143 VGND.n142 0.0565916
R756 uo_out[4] VGND.n491 0.0555
R757 VGND.n85 VGND.n84 0.0547113
R758 VGND.n100 VGND.n99 0.0546283
R759 VGND.n142 VGND.n140 0.0546283
R760 VGND.n456 VGND.n81 0.0545351
R761 VGND.n458 VGND.n457 0.0537058
R762 VGND.n378 VGND.n377 0.0505564
R763 VGND.n309 VGND.n308 0.0505564
R764 VGND.n102 VGND.n101 0.0497148
R765 VGND.n139 VGND.n138 0.0497148
R766 VGND.n84 VGND.n83 0.0483673
R767 VGND.n371 VGND.n102 0.0478846
R768 VGND.n138 VGND.n137 0.0478846
R769 VGND.n137 VGND.n136 0.04594
R770 VGND.n371 VGND.n370 0.04594
R771 VGND.n136 VGND.n135 0.0440235
R772 VGND.n370 VGND.n369 0.0440235
R773 VGND.n490 VGND.n1 0.043
R774 VGND.n446 VGND.n395 0.0425296
R775 VGND.n135 VGND.n134 0.0421344
R776 VGND.n369 VGND.n104 0.0421344
R777 VGND.n83 VGND.n82 0.0419304
R778 VGND.n176 VGND.n72 0.0411957
R779 VGND.n134 VGND.n133 0.0401312
R780 VGND.n365 VGND.n104 0.0401312
R781 VGND.n152 VGND.n151 0.0397586
R782 VGND.n389 VGND.n89 0.039235
R783 VGND.n133 VGND.n132 0.0386127
R784 VGND.n365 VGND.n364 0.0386127
R785 VGND.n132 VGND.n131 0.0365
R786 VGND.n364 VGND.n363 0.0365
R787 VGND.n462 VGND.n72 0.0356429
R788 VGND.n176 VGND.n175 0.0355141
R789 VGND.n131 VGND.n130 0.0351481
R790 VGND.n363 VGND.n106 0.0351481
R791 VGND.n175 VGND.n174 0.0337308
R792 VGND.n130 VGND.n129 0.0332724
R793 VGND.n359 VGND.n106 0.0332724
R794 VGND.n340 VGND.n339 0.032543
R795 VGND.n174 VGND.n173 0.0317753
R796 VGND.n129 VGND.n128 0.0313454
R797 VGND.n359 VGND.n358 0.0313454
R798 VGND.n351 VGND.n110 0.0307408
R799 VGND.n173 VGND.n172 0.0302379
R800 VGND.n128 VGND.n127 0.0299334
R801 VGND.n358 VGND.n357 0.0299334
R802 VGND.n324 VGND.n323 0.0298333
R803 VGND.n172 VGND.n171 0.0283213
R804 VGND.n127 VGND.n126 0.0279441
R805 VGND.n357 VGND.n108 0.0279441
R806 VGND.n80 VGND.n79 0.0273067
R807 VGND.n171 VGND.n170 0.0266297
R808 VGND.n126 VGND.n124 0.0263649
R809 VGND.n353 VGND.n108 0.0263649
R810 VGND.n170 VGND.n169 0.024961
R811 VGND.n443 VGND.n396 0.0249162
R812 VGND.n432 VGND.n425 0.0249162
R813 VGND.n124 VGND.n123 0.0247963
R814 VGND.n353 VGND.n352 0.0247963
R815 VGND.n169 VGND.n168 0.0233919
R816 VGND.n375 VGND.n372 0.02322
R817 VGND.n123 VGND.n122 0.0231622
R818 VGND.n352 VGND.n351 0.0231622
R819 VGND.n168 VGND.n167 0.0218333
R820 VGND.n246 VGND.n230 0.02175
R821 VGND.n27 VGND.n13 0.02175
R822 VGND.n58 VGND.n57 0.02175
R823 VGND.n445 VGND.n444 0.02162
R824 VGND.n426 VGND.n86 0.02162
R825 VGND.n122 VGND.n121 0.02162
R826 VGND.n462 VGND.n461 0.0212439
R827 VGND.n296 VGND.n295 0.0200345
R828 VGND.n167 VGND.n166 0.0199247
R829 VGND.n121 VGND.n120 0.0197957
R830 VGND.n166 VGND.n165 0.0186867
R831 VGND.n120 VGND.n119 0.0185662
R832 VGND.n457 VGND.n456 0.0170759
R833 VGND.n190 VGND.n165 0.0168721
R834 VGND.n119 VGND.n118 0.016764
R835 VGND.n0 uo_out[5] 0.0157601
R836 VGND.n400 uo_out[6] 0.0157601
R837 VGND.n401 uo_out[7] 0.0157601
R838 VGND.n402 uio_out[0] 0.0157601
R839 VGND.n403 uio_out[1] 0.0157601
R840 VGND.n407 uio_out[2] 0.0157601
R841 VGND.n408 uio_out[3] 0.0157601
R842 VGND.n409 uio_out[4] 0.0157601
R843 VGND.n410 uio_out[5] 0.0157601
R844 VGND.n411 uio_out[6] 0.0157601
R845 VGND.n412 uio_out[7] 0.0157601
R846 VGND.n413 uio_oe[0] 0.0157601
R847 VGND.n414 uio_oe[1] 0.0157601
R848 VGND.n415 uio_oe[2] 0.0157601
R849 VGND.n416 uio_oe[3] 0.0157601
R850 VGND.n417 uio_oe[4] 0.0157601
R851 VGND.n418 uio_oe[5] 0.0157601
R852 VGND.n419 uio_oe[6] 0.0157601
R853 VGND.n420 uio_oe[7] 0.0157601
R854 VGND.n79 VGND.n78 0.0153179
R855 VGND.n191 VGND.n190 0.0150695
R856 VGND.n118 VGND.n117 0.0149737
R857 VGND.n117 VGND.n116 0.0138158
R858 uo_out[5] VGND.n0 0.0137
R859 uo_out[6] VGND.n400 0.0137
R860 uo_out[7] VGND.n401 0.0137
R861 uio_out[0] VGND.n402 0.0137
R862 uio_out[1] VGND.n403 0.0137
R863 uio_out[2] VGND.n407 0.0137
R864 uio_out[3] VGND.n408 0.0137
R865 uio_out[4] VGND.n409 0.0137
R866 uio_out[5] VGND.n410 0.0137
R867 uio_out[6] VGND.n411 0.0137
R868 uio_out[7] VGND.n412 0.0137
R869 uio_oe[0] VGND.n413 0.0137
R870 uio_oe[1] VGND.n414 0.0137
R871 uio_oe[2] VGND.n415 0.0137
R872 uio_oe[3] VGND.n416 0.0137
R873 uio_oe[4] VGND.n417 0.0137
R874 uio_oe[5] VGND.n418 0.0137
R875 uio_oe[6] VGND.n419 0.0137
R876 uio_oe[7] VGND.n420 0.0137
R877 VGND.n323 VGND.n322 0.0132838
R878 VGND.n441 VGND.n397 0.0131992
R879 VGND.n435 VGND.n427 0.0131992
R880 VGND.n443 VGND.n398 0.0131916
R881 VGND.n428 VGND.n425 0.0131916
R882 VGND.n428 VGND.n423 0.0131916
R883 VGND.n421 VGND.n398 0.0131916
R884 VGND.n421 VGND.n397 0.0130858
R885 VGND.n427 VGND.n423 0.0130858
R886 VGND.n82 VGND.n81 0.0121797
R887 VGND.n116 VGND.n115 0.012041
R888 VGND.n442 VGND.n422 0.0115476
R889 VGND.n439 VGND.n437 0.0115476
R890 VGND.n436 VGND.n424 0.0115476
R891 VGND.n433 VGND.n429 0.0115476
R892 VGND.n430 VGND.n424 0.0115476
R893 VGND.n434 VGND.n433 0.0115476
R894 VGND.n438 VGND.n422 0.0115476
R895 VGND.n440 VGND.n439 0.0115476
R896 VGND.n440 VGND.n399 0.0115476
R897 VGND.n434 VGND.n431 0.0115476
R898 VGND.n431 VGND.n430 0.0115476
R899 VGND.n438 VGND.n399 0.0115476
R900 VGND.n115 VGND.n114 0.0105654
R901 VGND.n405 VGND.n404 0.0105
R902 VGND.n459 VGND.n78 0.00934499
R903 VGND.n451 VGND.n450 0.00920833
R904 VGND.n114 VGND.n113 0.00883987
R905 VGND.n455 VGND.n82 0.00874622
R906 VGND.n454 VGND.n83 0.0077971
R907 VGND.n338 VGND.n113 0.00737948
R908 VGND.n453 VGND.n84 0.00643951
R909 VGND.n339 VGND.n338 0.00594625
R910 VGND.n191 VGND.n164 0.00588981
R911 VGND.n457 VGND.n80 0.00446192
R912 VGND.n452 VGND.n85 0.00434654
R913 VGND.n308 VGND.n307 0.00206612
R914 VGND.n238 VGND.n222 0.00166667
R915 VGND.n485 VGND.n7 0.00166667
R916 VGND.n49 VGND.n39 0.00166667
R917 VGND.t86 VGND.n238 0.00133332
R918 VGND.n485 VGND.t99 0.00133332
R919 VGND.n479 VGND.n49 0.00133332
R920 VGND.n220 VGND.n211 0.001
R921 VGND.n235 VGND.n220 0.001
R922 VGND.n236 VGND.n221 0.001
R923 VGND.n488 VGND.n3 0.001
R924 VGND.n488 VGND.n487 0.001
R925 VGND.n6 VGND.n4 0.001
R926 VGND.n37 VGND.n8 0.001
R927 VGND.n50 VGND.n37 0.001
R928 VGND.n51 VGND.n38 0.001
R929 VGND.t103 VGND.n211 0.001
R930 VGND.n235 VGND.n221 0.001
R931 VGND.n236 VGND.n222 0.001
R932 VGND.t86 VGND.n3 0.001
R933 VGND.n487 VGND.n4 0.001
R934 VGND.n7 VGND.n6 0.001
R935 VGND.t99 VGND.n8 0.001
R936 VGND.n50 VGND.n38 0.001
R937 VGND.n51 VGND.n39 0.001
R938 uo_out[1].n3 uo_out[1].t2 15.0005
R939 uo_out[1] uo_out[1].n3 13.4668
R940 uo_out[1].n2 uo_out[1].n1 9.01747
R941 uo_out[1].n2 uo_out[1] 8.9065
R942 uo_out[1].n0 uo_out[1].t0 8.53421
R943 uo_out[1].n0 uo_out[1].t1 6.13626
R944 uo_out[1].n1 uo_out[1].n0 0.100612
R945 uo_out[1].n1 uo_out[1] 0.0585899
R946 uo_out[1].n3 uo_out[1] 0.04098
R947 uo_out[1] uo_out[1].n2 0.00678571
R948 VDPWR.n11 VDPWR.t48 34.1026
R949 VDPWR.n9 VDPWR.t28 34.1026
R950 VDPWR.n3 VDPWR.t9 34.1026
R951 VDPWR.n103 VDPWR.t3 34.1026
R952 VDPWR.n102 VDPWR.t79 34.1026
R953 VDPWR.n100 VDPWR.t61 34.1026
R954 VDPWR.n99 VDPWR.t59 34.1026
R955 VDPWR.n58 VDPWR.t76 34.1026
R956 VDPWR.n156 VDPWR.t5 34.1026
R957 VDPWR.n35 VDPWR.t32 34.1026
R958 VDPWR.n28 VDPWR.t0 34.1026
R959 VDPWR.n191 VDPWR.t55 34.1026
R960 VDPWR.n204 VDPWR.t35 34.1026
R961 VDPWR.n202 VDPWR.t81 34.1026
R962 VDPWR.n77 VDPWR.t88 34.1026
R963 VDPWR.n98 VDPWR.t41 34.1026
R964 VDPWR.n101 VDPWR.t43 34.1026
R965 VDPWR.n104 VDPWR.t22 34.1026
R966 VDPWR.n105 VDPWR.t30 34.1026
R967 VDPWR.n1 VDPWR.t7 34.1026
R968 VDPWR.n0 VDPWR.t24 34.1026
R969 VDPWR.n271 VDPWR.n214 19.7403
R970 VDPWR VDPWR.n11 18.2059
R971 VDPWR VDPWR.n9 18.2059
R972 VDPWR VDPWR.n3 18.2059
R973 VDPWR VDPWR.n103 18.2059
R974 VDPWR VDPWR.n102 18.2059
R975 VDPWR VDPWR.n100 18.2059
R976 VDPWR VDPWR.n99 18.2059
R977 VDPWR VDPWR.n58 18.2059
R978 VDPWR VDPWR.n156 18.2059
R979 VDPWR VDPWR.n35 18.2059
R980 VDPWR VDPWR.n28 18.2059
R981 VDPWR VDPWR.n191 18.2059
R982 VDPWR VDPWR.n204 18.2059
R983 VDPWR VDPWR.n202 18.2059
R984 VDPWR VDPWR.n77 18.2059
R985 VDPWR VDPWR.n98 18.2059
R986 VDPWR VDPWR.n101 18.2059
R987 VDPWR VDPWR.n104 18.2059
R988 VDPWR VDPWR.n105 18.2059
R989 VDPWR VDPWR.n1 18.2059
R990 VDPWR VDPWR.n0 18.2059
R991 VDPWR.n271 VDPWR.n270 18.0005
R992 VDPWR.n261 VDPWR.t34 17.378
R993 VDPWR.n248 VDPWR.t40 17.378
R994 VDPWR.n231 VDPWR.t45 17.378
R995 VDPWR.n262 VDPWR.t15 17.3693
R996 VDPWR.n246 VDPWR.t19 17.3693
R997 VDPWR.n230 VDPWR.t13 17.3693
R998 VDPWR.n11 VDPWR.t49 17.0233
R999 VDPWR.n9 VDPWR.t29 17.0233
R1000 VDPWR.n3 VDPWR.t10 17.0233
R1001 VDPWR.n103 VDPWR.t4 17.0233
R1002 VDPWR.n102 VDPWR.t80 17.0233
R1003 VDPWR.n100 VDPWR.t62 17.0233
R1004 VDPWR.n99 VDPWR.t60 17.0233
R1005 VDPWR.n58 VDPWR.t77 17.0233
R1006 VDPWR.n156 VDPWR.t6 17.0233
R1007 VDPWR.n35 VDPWR.t33 17.0233
R1008 VDPWR.n28 VDPWR.t1 17.0233
R1009 VDPWR.n191 VDPWR.t56 17.0233
R1010 VDPWR.n204 VDPWR.t36 17.0233
R1011 VDPWR.n202 VDPWR.t82 17.0233
R1012 VDPWR.n77 VDPWR.t89 17.0233
R1013 VDPWR.n98 VDPWR.t42 17.0233
R1014 VDPWR.n101 VDPWR.t44 17.0233
R1015 VDPWR.n104 VDPWR.t23 17.0233
R1016 VDPWR.n105 VDPWR.t31 17.0233
R1017 VDPWR.n1 VDPWR.t8 17.0233
R1018 VDPWR.n0 VDPWR.t25 17.0233
R1019 VDPWR.n261 VDPWR.t18 17.0005
R1020 VDPWR.t12 VDPWR.n229 17.0005
R1021 VDPWR.n268 VDPWR.t12 17.0005
R1022 VDPWR.n248 VDPWR.t14 17.0005
R1023 VDPWR.t11 VDPWR.n250 17.0005
R1024 VDPWR.t11 VDPWR.n252 17.0005
R1025 VDPWR.t11 VDPWR.n241 17.0005
R1026 VDPWR.n231 VDPWR.t20 17.0005
R1027 VDPWR.t12 VDPWR.n215 17.0005
R1028 VDPWR.t12 VDPWR.n222 17.0005
R1029 VDPWR.t12 VDPWR.n235 17.0005
R1030 VDPWR.n264 VDPWR.t11 17.0005
R1031 VDPWR.n272 VDPWR.n271 12.4694
R1032 VDPWR.n212 VDPWR.n211 9.2117
R1033 VDPWR.n208 VDPWR.n194 9.18823
R1034 VDPWR.n212 VDPWR.n22 9.18823
R1035 VDPWR.n212 VDPWR.n21 9.05079
R1036 VDPWR.n209 VDPWR.n208 9.0005
R1037 VDPWR.n210 VDPWR.n22 9.0005
R1038 VDPWR.n209 VDPWR.n25 9.0005
R1039 VDPWR.n210 VDPWR.n21 9.0005
R1040 VDPWR.n209 VDPWR.n23 9.0005
R1041 VDPWR.n211 VDPWR.n210 9.0005
R1042 VDPWR.n199 VDPWR.n198 9.0005
R1043 VDPWR.n196 VDPWR.n15 9.0005
R1044 VDPWR.n276 VDPWR.n17 9.0005
R1045 VDPWR.n259 VDPWR.t65 8.80285
R1046 VDPWR.n237 VDPWR.t69 8.80285
R1047 VDPWR.n225 VDPWR.t52 8.80285
R1048 VDPWR.t2 VDPWR.n242 8.501
R1049 VDPWR.t11 VDPWR.n256 8.47111
R1050 VDPWR.t11 VDPWR.n258 8.47111
R1051 VDPWR.t12 VDPWR.n226 8.47111
R1052 VDPWR.t12 VDPWR.n219 8.47111
R1053 VDPWR.t12 VDPWR.n217 8.47111
R1054 VDPWR.n266 VDPWR.n238 8.47111
R1055 VDPWR.n265 VDPWR.n239 8.47111
R1056 VDPWR.n224 VDPWR.t50 6.07323
R1057 VDPWR.n257 VDPWR.t63 6.073
R1058 VDPWR.n218 VDPWR.t68 6.073
R1059 VDPWR.n107 VDPWR.n106 6.01045
R1060 VDPWR.n228 VDPWR.t38 5.98925
R1061 VDPWR.n216 VDPWR.t37 5.98882
R1062 VDPWR.n255 VDPWR.t86 5.98825
R1063 VDPWR.n253 VDPWR.t85 5.98825
R1064 VDPWR.n220 VDPWR.t46 5.98825
R1065 VDPWR.n234 VDPWR.t47 5.98825
R1066 VDPWR.n109 VDPWR.n108 5.98145
R1067 VDPWR.n10 VDPWR 5.96901
R1068 VDPWR.n192 VDPWR.n190 5.84778
R1069 VDPWR.t12 VDPWR.n227 5.61485
R1070 VDPWR.t11 VDPWR.n254 5.61485
R1071 VDPWR.t12 VDPWR.n221 5.61485
R1072 VDPWR.t12 VDPWR.n267 5.61485
R1073 VDPWR.n273 VDPWR 5.2541
R1074 VDPWR.n112 VDPWR.n111 5.21746
R1075 VDPWR.n4 VDPWR 4.89941
R1076 VDPWR.n280 VDPWR 4.6152
R1077 VDPWR.n194 VDPWR.n193 4.53071
R1078 VDPWR.n207 VDPWR.n26 4.51901
R1079 VDPWR.n206 VDPWR.n20 4.50989
R1080 VDPWR VDPWR.n291 4.13588
R1081 VDPWR.n2 VDPWR 3.92388
R1082 VDPWR.n107 VDPWR 3.88095
R1083 VDPWR.n106 VDPWR 3.84419
R1084 VDPWR.n203 VDPWR 3.78722
R1085 VDPWR.n108 VDPWR 3.41222
R1086 VDPWR.t11 VDPWR.n251 3.33162
R1087 VDPWR.t12 VDPWR.n233 3.30723
R1088 VDPWR.t11 VDPWR.n247 3.30706
R1089 VDPWR.n205 VDPWR 3.28289
R1090 VDPWR.n198 VDPWR.n197 3.0005
R1091 VDPWR.n15 VDPWR.n13 3.0005
R1092 VDPWR.n277 VDPWR.n276 3.0005
R1093 VDPWR.n192 VDPWR 2.98934
R1094 VDPWR.t11 VDPWR.n263 2.72512
R1095 VDPWR.n280 VDPWR.n279 2.5318
R1096 VDPWR.n29 VDPWR 2.53128
R1097 VDPWR.n155 VDPWR.n57 2.46388
R1098 VDPWR.n109 VDPWR 2.33518
R1099 VDPWR.t11 VDPWR.n245 2.29759
R1100 VDPWR.n194 VDPWR.n24 2.27162
R1101 VDPWR.n195 VDPWR.n16 2.26628
R1102 VDPWR.n213 VDPWR.n212 2.2505
R1103 VDPWR.n209 VDPWR.n24 2.2505
R1104 VDPWR.n210 VDPWR.n19 2.2505
R1105 VDPWR.n274 VDPWR.n16 2.2505
R1106 VDPWR.n276 VDPWR.n275 2.2505
R1107 VDPWR.n244 VDPWR 2.0605
R1108 VDPWR.n36 VDPWR 1.94477
R1109 VDPWR.n273 VDPWR.n272 1.89976
R1110 VDPWR.n110 VDPWR 1.74056
R1111 VDPWR.n112 VDPWR 1.53994
R1112 VDPWR.n240 VDPWR 1.53643
R1113 VDPWR.n274 VDPWR.n273 1.47736
R1114 VDPWR.n272 VDPWR.n213 1.46416
R1115 VDPWR.n111 VDPWR 1.39911
R1116 VDPWR.n157 VDPWR 1.30374
R1117 VDPWR.n114 VDPWR 1.19117
R1118 VDPWR.n275 VDPWR.n18 1.14638
R1119 VDPWR.n113 VDPWR.n112 0.923201
R1120 VDPWR.n135 VDPWR 0.895684
R1121 VDPWR.n154 VDPWR 0.886
R1122 VDPWR.n225 VDPWR.n223 0.854038
R1123 VDPWR.n260 VDPWR.n259 0.851125
R1124 VDPWR.n262 VDPWR.n260 0.805789
R1125 VDPWR.n230 VDPWR.n223 0.803932
R1126 VDPWR.t12 VDPWR.n223 0.802654
R1127 VDPWR.t11 VDPWR.n260 0.800901
R1128 VDPWR.n291 VDPWR.n290 0.762687
R1129 VDPWR.n269 VDPWR 0.543
R1130 VDPWR.n185 VDPWR.n27 0.531002
R1131 VDPWR.n169 VDPWR.n168 0.507992
R1132 VDPWR.n84 VDPWR.n83 0.507992
R1133 VDPWR.n263 VDPWR.n261 0.410237
R1134 VDPWR.n110 VDPWR.n109 0.409089
R1135 VDPWR.t2 VDPWR.n236 0.40574
R1136 VDPWR.n245 VDPWR.n244 0.392162
R1137 VDPWR.n263 VDPWR.n262 0.389189
R1138 VDPWR.n246 VDPWR.n245 0.374189
R1139 VDPWR.n106 VDPWR.n2 0.363276
R1140 VDPWR.n205 VDPWR.n203 0.348974
R1141 VDPWR.n243 VDPWR.t2 0.341
R1142 VDPWR.n233 VDPWR.n230 0.336433
R1143 VDPWR.n247 VDPWR.n246 0.336118
R1144 VDPWR.n111 VDPWR.n110 0.332665
R1145 VDPWR.n249 VDPWR.n247 0.331746
R1146 VDPWR.n233 VDPWR.n232 0.331445
R1147 VDPWR.n59 VDPWR.n57 0.330588
R1148 VDPWR.n108 VDPWR.n107 0.323555
R1149 VDPWR.n158 VDPWR.n155 0.313098
R1150 VDPWR.n206 VDPWR.n205 0.312824
R1151 VDPWR.n267 VDPWR.n266 0.300775
R1152 VDPWR.n291 VDPWR.n2 0.289257
R1153 VDPWR.n170 VDPWR.n169 0.2887
R1154 VDPWR.n85 VDPWR.n84 0.2887
R1155 VDPWR.n60 VDPWR.n59 0.280623
R1156 VDPWR.n251 VDPWR 0.273551
R1157 VDPWR.n184 VDPWR.n30 0.251853
R1158 VDPWR.n183 VDPWR.n31 0.2469
R1159 VDPWR.n182 VDPWR.n32 0.24161
R1160 VDPWR.n115 VDPWR.n97 0.24161
R1161 VDPWR.n266 VDPWR.n265 0.241078
R1162 VDPWR.n61 VDPWR.n60 0.240286
R1163 VDPWR.n181 VDPWR.n33 0.237849
R1164 VDPWR.n116 VDPWR.n96 0.237849
R1165 VDPWR.n180 VDPWR.n34 0.234669
R1166 VDPWR.n117 VDPWR.n95 0.234669
R1167 VDPWR.n179 VDPWR.n36 0.231561
R1168 VDPWR.n118 VDPWR.n94 0.231561
R1169 VDPWR.n189 VDPWR.n188 0.230306
R1170 VDPWR.n178 VDPWR.n37 0.226786
R1171 VDPWR.n119 VDPWR.n93 0.226786
R1172 VDPWR.n171 VDPWR.n170 0.225081
R1173 VDPWR.n86 VDPWR.n85 0.225081
R1174 VDPWR.n177 VDPWR.n38 0.22337
R1175 VDPWR.n120 VDPWR.n92 0.22337
R1176 VDPWR.n176 VDPWR.n39 0.219324
R1177 VDPWR.n121 VDPWR.n91 0.219324
R1178 VDPWR.n175 VDPWR.n40 0.217223
R1179 VDPWR.n122 VDPWR.n90 0.217223
R1180 VDPWR.n174 VDPWR.n41 0.213359
R1181 VDPWR.n123 VDPWR.n89 0.213359
R1182 VDPWR.n186 VDPWR.n185 0.212767
R1183 VDPWR.n211 VDPWR.n23 0.2117
R1184 VDPWR.n173 VDPWR.n42 0.211333
R1185 VDPWR.n124 VDPWR.n88 0.211333
R1186 VDPWR.n172 VDPWR.n43 0.208253
R1187 VDPWR.n125 VDPWR.n87 0.208253
R1188 VDPWR VDPWR.n251 0.205841
R1189 VDPWR.n62 VDPWR.n61 0.204702
R1190 VDPWR.n171 VDPWR.n44 0.204642
R1191 VDPWR.n126 VDPWR.n86 0.204642
R1192 VDPWR.n170 VDPWR.n45 0.202722
R1193 VDPWR.n127 VDPWR.n85 0.202722
R1194 VDPWR.n190 VDPWR.n27 0.201278
R1195 VDPWR.n169 VDPWR.n46 0.19982
R1196 VDPWR.n128 VDPWR.n84 0.19982
R1197 VDPWR.n159 VDPWR.n158 0.193685
R1198 VDPWR.n63 VDPWR.n62 0.187779
R1199 VDPWR.n267 VDPWR.n237 0.185825
R1200 VDPWR.n265 VDPWR.n264 0.180789
R1201 VDPWR.n172 VDPWR.n171 0.177266
R1202 VDPWR.n87 VDPWR.n86 0.177266
R1203 VDPWR.n64 VDPWR.n63 0.175509
R1204 VDPWR.n167 VDPWR.n48 0.173049
R1205 VDPWR.n130 VDPWR.n82 0.173049
R1206 VDPWR.n166 VDPWR.n49 0.172207
R1207 VDPWR.n131 VDPWR.n81 0.172207
R1208 VDPWR.n256 VDPWR.n255 0.172039
R1209 VDPWR.n220 VDPWR.n219 0.172039
R1210 VDPWR.n165 VDPWR.n50 0.171374
R1211 VDPWR.n132 VDPWR.n80 0.171374
R1212 VDPWR.n164 VDPWR.n51 0.169731
R1213 VDPWR.n133 VDPWR.n79 0.169731
R1214 VDPWR.n163 VDPWR.n52 0.168921
R1215 VDPWR.n134 VDPWR.n78 0.168921
R1216 VDPWR.n201 VDPWR.n200 0.168402
R1217 VDPWR.n162 VDPWR.n53 0.167325
R1218 VDPWR.n135 VDPWR.n76 0.167325
R1219 VDPWR.n290 VDPWR.n289 0.166596
R1220 VDPWR.n161 VDPWR.n54 0.166538
R1221 VDPWR.n136 VDPWR.n75 0.166538
R1222 VDPWR.n160 VDPWR.n55 0.165758
R1223 VDPWR.n137 VDPWR.n74 0.165758
R1224 VDPWR.n113 VDPWR.n97 0.165337
R1225 VDPWR.n159 VDPWR.n56 0.164986
R1226 VDPWR.n138 VDPWR.n73 0.164986
R1227 VDPWR.n139 VDPWR.n72 0.164221
R1228 VDPWR.n140 VDPWR.n71 0.163463
R1229 VDPWR.n188 VDPWR.n187 0.162204
R1230 VDPWR.n142 VDPWR.n69 0.161968
R1231 VDPWR.n141 VDPWR.n70 0.161968
R1232 VDPWR.n144 VDPWR.n67 0.161231
R1233 VDPWR.n143 VDPWR.n68 0.161231
R1234 VDPWR.n147 VDPWR.n64 0.159776
R1235 VDPWR.n146 VDPWR.n65 0.159776
R1236 VDPWR.n145 VDPWR.n66 0.159776
R1237 VDPWR.n149 VDPWR.n62 0.159059
R1238 VDPWR.n148 VDPWR.n63 0.159059
R1239 VDPWR.n152 VDPWR.n59 0.158348
R1240 VDPWR.n151 VDPWR.n60 0.158348
R1241 VDPWR.n150 VDPWR.n61 0.158348
R1242 VDPWR.n65 VDPWR.n64 0.157911
R1243 VDPWR.n173 VDPWR.n172 0.157621
R1244 VDPWR.n88 VDPWR.n87 0.157621
R1245 VDPWR.n153 VDPWR.n57 0.154546
R1246 VDPWR.n168 VDPWR.n47 0.15242
R1247 VDPWR.n129 VDPWR.n83 0.15242
R1248 VDPWR.n282 VDPWR.n281 0.152188
R1249 VDPWR.n66 VDPWR.n65 0.147308
R1250 VDPWR.n207 VDPWR.n22 0.147167
R1251 VDPWR.n67 VDPWR.n66 0.14126
R1252 VDPWR.n174 VDPWR.n173 0.141098
R1253 VDPWR.n89 VDPWR.n88 0.141098
R1254 VDPWR.n258 VDPWR.n257 0.140789
R1255 VDPWR.n218 VDPWR.n217 0.140789
R1256 VDPWR.n226 VDPWR.n224 0.140789
R1257 VDPWR.n290 VDPWR.n4 0.137615
R1258 VDPWR.n249 VDPWR.n248 0.136382
R1259 VDPWR.n232 VDPWR.n231 0.136382
R1260 VDPWR.n287 VDPWR.n5 0.135022
R1261 VDPWR.n68 VDPWR.n67 0.133682
R1262 VDPWR.n227 VDPWR.n216 0.129236
R1263 VDPWR.n255 VDPWR.n254 0.129236
R1264 VDPWR.n221 VDPWR.n220 0.129236
R1265 VDPWR.n228 VDPWR.n227 0.128325
R1266 VDPWR.n254 VDPWR.n253 0.128325
R1267 VDPWR.n234 VDPWR.n221 0.128325
R1268 VDPWR.n69 VDPWR.n68 0.127233
R1269 VDPWR.n186 VDPWR.n30 0.1269
R1270 VDPWR.n175 VDPWR.n174 0.126475
R1271 VDPWR.n90 VDPWR.n89 0.126475
R1272 VDPWR.n70 VDPWR.n69 0.123269
R1273 VDPWR.n71 VDPWR.n70 0.121562
R1274 VDPWR.n193 VDPWR.n23 0.1171
R1275 VDPWR.n72 VDPWR.n71 0.116891
R1276 VDPWR.n176 VDPWR.n175 0.116337
R1277 VDPWR.n91 VDPWR.n90 0.116337
R1278 VDPWR.n259 VDPWR.n258 0.115789
R1279 VDPWR.n237 VDPWR.n217 0.115789
R1280 VDPWR.n226 VDPWR.n225 0.115789
R1281 VDPWR.n73 VDPWR.n72 0.114401
R1282 VDPWR.n229 VDPWR.n228 0.113
R1283 VDPWR.n253 VDPWR.n252 0.113
R1284 VDPWR.n235 VDPWR.n234 0.113
R1285 VDPWR.n268 VDPWR.n216 0.11175
R1286 VDPWR.n160 VDPWR.n159 0.111106
R1287 VDPWR.n74 VDPWR.n73 0.111106
R1288 VDPWR.n161 VDPWR.n160 0.110556
R1289 VDPWR.n75 VDPWR.n74 0.110556
R1290 VDPWR.n162 VDPWR.n161 0.108981
R1291 VDPWR.n76 VDPWR.n75 0.108981
R1292 VDPWR.n78 VDPWR.n76 0.108669
R1293 VDPWR.n79 VDPWR.n78 0.108583
R1294 VDPWR.n177 VDPWR.n176 0.108277
R1295 VDPWR.n92 VDPWR.n91 0.108277
R1296 VDPWR.n80 VDPWR.n79 0.108072
R1297 VDPWR.n163 VDPWR.n162 0.107646
R1298 VDPWR.n164 VDPWR.n163 0.107594
R1299 VDPWR.n82 VDPWR.n81 0.107345
R1300 VDPWR.n166 VDPWR.n165 0.107234
R1301 VDPWR.n81 VDPWR.n80 0.107234
R1302 VDPWR.n165 VDPWR.n164 0.107115
R1303 VDPWR.n167 VDPWR.n166 0.106465
R1304 VDPWR.n178 VDPWR.n177 0.103826
R1305 VDPWR.n93 VDPWR.n92 0.103826
R1306 VDPWR.n257 VDPWR.n256 0.100789
R1307 VDPWR.n219 VDPWR.n218 0.100789
R1308 VDPWR.n179 VDPWR.n178 0.0994295
R1309 VDPWR.n94 VDPWR.n93 0.0994295
R1310 VDPWR.n180 VDPWR.n179 0.096586
R1311 VDPWR.n95 VDPWR.n94 0.096586
R1312 VDPWR.n284 VDPWR.n8 0.0942964
R1313 VDPWR.n181 VDPWR.n180 0.0929227
R1314 VDPWR.n96 VDPWR.n95 0.0929227
R1315 VDPWR.n182 VDPWR.n181 0.0912154
R1316 VDPWR.n97 VDPWR.n96 0.0912154
R1317 VDPWR.n6 VDPWR.n5 0.0893224
R1318 VDPWR.n183 VDPWR.n182 0.0884738
R1319 VDPWR.n270 VDPWR.n269 0.088
R1320 VDPWR.n184 VDPWR.n183 0.0871337
R1321 VDPWR.n185 VDPWR.n184 0.0864426
R1322 VDPWR.n31 VDPWR.n30 0.0816497
R1323 VDPWR.n187 VDPWR.n186 0.0787288
R1324 VDPWR.n32 VDPWR.n31 0.0781471
R1325 VDPWR.n115 VDPWR.n114 0.0781471
R1326 VDPWR.n288 VDPWR.n287 0.0761377
R1327 VDPWR.n33 VDPWR.n32 0.0757832
R1328 VDPWR.n116 VDPWR.n115 0.0757832
R1329 VDPWR.n34 VDPWR.n33 0.0734143
R1330 VDPWR.n117 VDPWR.n116 0.0734143
R1331 VDPWR.n287 VDPWR.n286 0.0722058
R1332 VDPWR.n240 VDPWR.n214 0.0717963
R1333 VDPWR.n283 VDPWR.n10 0.071653
R1334 VDPWR.n36 VDPWR.n34 0.071596
R1335 VDPWR.n118 VDPWR.n117 0.071596
R1336 VDPWR.n37 VDPWR.n36 0.0688352
R1337 VDPWR.n119 VDPWR.n118 0.0688352
R1338 VDPWR.n48 VDPWR.n47 0.0683607
R1339 VDPWR.n130 VDPWR.n129 0.0683607
R1340 VDPWR.n284 VDPWR.n283 0.0679195
R1341 VDPWR.n38 VDPWR.n37 0.0662582
R1342 VDPWR.n120 VDPWR.n119 0.0662582
R1343 VDPWR.n244 VDPWR.n241 0.0656852
R1344 VDPWR.n188 VDPWR.n27 0.0656852
R1345 VDPWR.n39 VDPWR.n38 0.0641087
R1346 VDPWR.n121 VDPWR.n120 0.0641087
R1347 VDPWR.n114 VDPWR.n113 0.0637952
R1348 VDPWR.n197 VDPWR.n12 0.0627642
R1349 VDPWR.n200 VDPWR.n199 0.0624718
R1350 VDPWR.n40 VDPWR.n39 0.0612059
R1351 VDPWR.n122 VDPWR.n121 0.0612059
R1352 VDPWR.n229 VDPWR 0.0605
R1353 VDPWR.n252 VDPWR 0.0605
R1354 VDPWR VDPWR.n250 0.0605
R1355 VDPWR.n235 VDPWR 0.0605
R1356 VDPWR VDPWR.n222 0.0605
R1357 VDPWR.n41 VDPWR.n40 0.0599468
R1358 VDPWR.n123 VDPWR.n122 0.0599468
R1359 VDPWR.n285 VDPWR.n7 0.0577377
R1360 VDPWR.n42 VDPWR.n41 0.0571702
R1361 VDPWR.n124 VDPWR.n123 0.0571702
R1362 VDPWR.n43 VDPWR.n42 0.0555
R1363 VDPWR.n125 VDPWR.n124 0.0555
R1364 VDPWR.n44 VDPWR.n43 0.0535722
R1365 VDPWR.n126 VDPWR.n125 0.0535722
R1366 VDPWR.n281 VDPWR.n280 0.0532395
R1367 VDPWR.n288 VDPWR.n4 0.0528027
R1368 VDPWR.n289 VDPWR.n288 0.0522
R1369 VDPWR.n45 VDPWR.n44 0.0509772
R1370 VDPWR.n127 VDPWR.n126 0.0509772
R1371 VDPWR.n46 VDPWR.n45 0.0493889
R1372 VDPWR.n128 VDPWR.n127 0.0493889
R1373 VDPWR.n47 VDPWR.n46 0.04758
R1374 VDPWR.n129 VDPWR.n128 0.04758
R1375 VDPWR.n279 VDPWR.n12 0.0460752
R1376 VDPWR.n190 VDPWR.n189 0.045577
R1377 VDPWR.n168 VDPWR.n167 0.0448348
R1378 VDPWR.n83 VDPWR.n82 0.0448348
R1379 VDPWR.n49 VDPWR.n48 0.0427745
R1380 VDPWR.n131 VDPWR.n130 0.0427745
R1381 VDPWR.n283 VDPWR.n282 0.0419028
R1382 VDPWR.n208 VDPWR.n207 0.0415667
R1383 VDPWR.n200 VDPWR.n12 0.0413571
R1384 VDPWR.n285 VDPWR.n284 0.0410333
R1385 VDPWR.n279 VDPWR.n278 0.0408577
R1386 VDPWR.n50 VDPWR.n49 0.0408512
R1387 VDPWR.n132 VDPWR.n131 0.0408512
R1388 VDPWR.n224 VDPWR.n215 0.0405
R1389 VDPWR.n197 VDPWR.n13 0.0403491
R1390 VDPWR.n199 VDPWR.n196 0.040162
R1391 VDPWR.n196 VDPWR.n17 0.040162
R1392 VDPWR.n207 VDPWR.n21 0.0397857
R1393 VDPWR.n51 VDPWR.n50 0.0389466
R1394 VDPWR.n133 VDPWR.n132 0.0389466
R1395 VDPWR.n207 VDPWR.n206 0.0385976
R1396 VDPWR.n187 VDPWR.n29 0.0383925
R1397 VDPWR.n52 VDPWR.n51 0.0377308
R1398 VDPWR.n134 VDPWR.n133 0.0377308
R1399 VDPWR.n189 VDPWR.n29 0.0376329
R1400 VDPWR.n53 VDPWR.n52 0.0358684
R1401 VDPWR.n135 VDPWR.n134 0.0358684
R1402 VDPWR.n286 VDPWR.n285 0.0356133
R1403 VDPWR.n278 VDPWR.n13 0.0341226
R1404 VDPWR.n54 VDPWR.n53 0.0338649
R1405 VDPWR.n136 VDPWR.n135 0.0338649
R1406 VDPWR.n55 VDPWR.n54 0.0320472
R1407 VDPWR.n137 VDPWR.n136 0.0320472
R1408 VDPWR.n56 VDPWR.n55 0.0306596
R1409 VDPWR.n138 VDPWR.n137 0.0306596
R1410 VDPWR.n270 VDPWR.n215 0.0305
R1411 VDPWR.n157 VDPWR.n56 0.0288738
R1412 VDPWR.n139 VDPWR.n138 0.0288738
R1413 VDPWR.n193 VDPWR.n25 0.0282619
R1414 VDPWR.n140 VDPWR.n139 0.0271047
R1415 VDPWR.n250 VDPWR.n249 0.02675
R1416 VDPWR.n232 VDPWR.n222 0.02675
R1417 VDPWR.n141 VDPWR.n140 0.0257593
R1418 VDPWR.n264 VDPWR.n240 0.0255
R1419 VDPWR.n210 VDPWR.n209 0.0249162
R1420 VDPWR.n276 VDPWR.n15 0.0249162
R1421 VDPWR.n276 VDPWR.n16 0.0249162
R1422 VDPWR.n142 VDPWR.n141 0.0239128
R1423 VDPWR.n155 VDPWR.n154 0.02261
R1424 VDPWR.n203 VDPWR.n201 0.0225381
R1425 VDPWR.n143 VDPWR.n142 0.0222982
R1426 VDPWR.n24 VDPWR.n19 0.02162
R1427 VDPWR.n213 VDPWR.n19 0.02162
R1428 VDPWR.n275 VDPWR.n274 0.02162
R1429 VDPWR.n144 VDPWR.n143 0.0205913
R1430 VDPWR.n145 VDPWR.n144 0.018984
R1431 VDPWR.n282 VDPWR.n8 0.0188236
R1432 VDPWR.n158 VDPWR.n157 0.018557
R1433 VDPWR.n193 VDPWR.n192 0.0182408
R1434 VDPWR.n154 VDPWR.n153 0.0179271
R1435 VDPWR.n146 VDPWR.n145 0.0176222
R1436 VDPWR.n201 VDPWR.n195 0.0170391
R1437 VDPWR.n147 VDPWR.n146 0.0160294
R1438 VDPWR.n289 VDPWR.n5 0.015852
R1439 VDPWR.n8 VDPWR.n7 0.0156247
R1440 VDPWR.n281 VDPWR.n10 0.0149236
R1441 VDPWR.n7 VDPWR.n6 0.0148367
R1442 VDPWR.n148 VDPWR.n147 0.0140385
R1443 VDPWR.n198 VDPWR.n18 0.0138871
R1444 VDPWR.n18 VDPWR.n15 0.0133938
R1445 VDPWR.n194 VDPWR.n26 0.0132264
R1446 VDPWR.n212 VDPWR.n20 0.0132264
R1447 VDPWR.n149 VDPWR.n148 0.0131847
R1448 VDPWR.n209 VDPWR.n26 0.0131568
R1449 VDPWR.n210 VDPWR.n20 0.0131568
R1450 VDPWR.n207 VDPWR.n25 0.0115
R1451 VDPWR.n150 VDPWR.n149 0.0112027
R1452 VDPWR.n277 VDPWR.n14 0.0100472
R1453 VDPWR.n17 VDPWR.n14 0.0100023
R1454 VDPWR.n151 VDPWR.n150 0.00957623
R1455 VDPWR.n152 VDPWR.n151 0.00839238
R1456 VDPWR.n278 VDPWR.n277 0.00672642
R1457 VDPWR.n241 VDPWR.n214 0.00661111
R1458 VDPWR.n153 VDPWR.n152 0.00641928
R1459 VDPWR.n195 VDPWR.n14 0.00463323
R1460 VDPWR.n269 VDPWR.n268 0.003
R1461 VDPWR.n238 VDPWR.n236 0.00197617
R1462 VDPWR.n286 VDPWR.n6 0.00108355
R1463 VDPWR.t12 VDPWR.n236 0.00102381
R1464 VDPWR.n243 VDPWR.n239 0.001
R1465 VDPWR.n242 VDPWR.n239 0.001
R1466 VDPWR.t11 VDPWR.n243 0.001
R1467 VDPWR.n242 VDPWR.n238 0.001
R1468 uo_out[2].n3 uo_out[2].t2 15.0005
R1469 uo_out[2] uo_out[2].n3 12.8496
R1470 uo_out[2].n2 uo_out[2] 12.5614
R1471 uo_out[2].n2 uo_out[2].n1 9.01936
R1472 uo_out[2].n0 uo_out[2].t1 8.53421
R1473 uo_out[2].n0 uo_out[2].t0 6.13626
R1474 uo_out[2].n1 uo_out[2].n0 0.0993764
R1475 uo_out[2].n1 uo_out[2] 0.0598258
R1476 uo_out[2] uo_out[2].n2 0.0388429
R1477 uo_out[2].n3 uo_out[2] 0.02525
R1478 uo_out[0].n4 uo_out[0].n3 33.1637
R1479 uo_out[0].n5 uo_out[0].t1 18.0455
R1480 uo_out[0] uo_out[0].t0 18.0125
R1481 uo_out[0].n1 uo_out[0].t3 15.0005
R1482 uo_out[0].n2 uo_out[0].n1 9.03505
R1483 uo_out[0].n3 uo_out[0].n2 6.7505
R1484 uo_out[0].n5 uo_out[0].n4 6.67645
R1485 uo_out[0].n4 uo_out[0].n0 4.90955
R1486 uo_out[0].n0 uo_out[0].t2 3.93974
R1487 uo_out[0].n3 uo_out[0] 1.35863
R1488 uo_out[0] uo_out[0].n5 0.0885
R1489 uo_out[0].n0 uo_out[0] 0.0446962
R1490 uo_out[0].n2 uo_out[0] 0.0401
R1491 uo_out[0].n1 uo_out[0] 0.02525
R1492 uo_out[3].n2 uo_out[3] 15.6957
R1493 uo_out[3].n2 uo_out[3].n1 9.0225
R1494 uo_out[3].n0 uo_out[3].t1 8.53421
R1495 uo_out[3].n0 uo_out[3].t0 6.13626
R1496 uo_out[3].n1 uo_out[3].n0 0.11668
R1497 uo_out[3].n1 uo_out[3] 0.0425225
R1498 uo_out[3] uo_out[3].n2 0.0357
C10 uo_out[0] VGND 11.2531f
C11 VDPWR VGND 0.10247p
.ends

