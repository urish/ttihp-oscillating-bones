magic
tech ihp-sg13g2
magscale 1 2
timestamp 1741277038
<< metal1 >>
rect 14979 44173 15226 44269
rect 15322 44173 15332 44269
rect 14961 43919 15227 43977
rect 9158 43628 9176 43724
rect 9272 43628 9524 43724
rect 15169 43511 15227 43919
rect 12120 43453 15227 43511
rect 8882 43220 10590 43332
rect 8882 43014 8994 43220
rect 8896 32168 8996 41646
rect 10478 41442 10590 43220
rect 12120 43028 12178 43453
rect 12092 41478 12204 41630
rect 12036 41442 12046 41478
rect 10478 41330 12046 41442
rect 12036 41298 12046 41330
rect 12234 41298 12244 41478
rect 1494 22582 1504 22882
rect 1804 22582 1814 22882
<< via1 >>
rect 15226 44173 15322 44269
rect 9176 43628 9272 43724
rect 12046 41298 12234 41478
rect 1504 22582 1804 22882
<< metal2 >>
rect 14044 44818 14108 44828
rect 14044 44728 14108 44738
rect 14596 44818 14660 44828
rect 14596 44728 14660 44738
rect 15148 44818 15212 44828
rect 14046 44554 14098 44728
rect 9738 44502 14098 44554
rect 9738 43760 9790 44502
rect 14600 44450 14652 44728
rect 11680 44398 14652 44450
rect 9152 43724 9312 43756
rect 11680 43752 11732 44398
rect 15148 44366 15212 44738
rect 13608 44314 15212 44366
rect 13608 43772 13660 44314
rect 15226 44269 15322 44279
rect 15226 44163 15322 44173
rect 14952 43980 15012 43990
rect 14952 43890 15012 43900
rect 9152 43628 9176 43724
rect 9272 43628 9312 43724
rect 9152 43584 9312 43628
rect 9152 43424 10629 43584
rect 7118 43026 7230 43036
rect 10469 43026 10629 43424
rect 13450 43352 13618 43362
rect 13448 43240 13450 43350
rect 13618 43240 13626 43350
rect 7230 42914 7632 43026
rect 10283 42936 10819 43026
rect 13448 42914 13626 43240
rect 7118 42904 7230 42914
rect 12046 41478 12234 41488
rect 12046 41288 12234 41298
rect 6372 23314 6672 23324
rect 6372 23004 6672 23014
rect 1504 22882 1804 22892
rect 1804 22582 2304 22882
rect 1504 22572 1804 22582
<< via2 >>
rect 14044 44738 14108 44818
rect 14596 44738 14660 44818
rect 15148 44738 15212 44818
rect 15226 44173 15322 44269
rect 14952 43900 15012 43980
rect 9176 43628 9272 43724
rect 13450 43240 13618 43352
rect 7118 42914 7230 43026
rect 12046 41298 12234 41478
rect 6372 23014 6672 23314
rect 1504 22582 1804 22882
<< metal3 >>
rect 14034 44818 14118 44853
rect 14034 44738 14044 44818
rect 14108 44738 14118 44818
rect 14034 44733 14118 44738
rect 14586 44818 14670 44853
rect 14586 44738 14596 44818
rect 14660 44738 14670 44818
rect 14586 44733 14670 44738
rect 15138 44818 15222 44853
rect 15138 44738 15148 44818
rect 15212 44738 15222 44818
rect 15138 44733 15222 44738
rect 15216 44272 15332 44274
rect 15184 44269 15384 44272
rect 15184 44173 15226 44269
rect 15322 44173 15384 44269
rect 14932 43980 15032 44000
rect 14932 43900 14950 43980
rect 15014 43900 15032 43980
rect 14932 43880 15032 43900
rect 9154 43729 9292 43746
rect 9154 43623 9171 43729
rect 9277 43623 9292 43729
rect 9154 43606 9292 43623
rect 15184 43410 15384 44173
rect 624 43408 15384 43410
rect 624 43210 658 43408
rect 648 43208 658 43210
rect 858 43352 15384 43408
rect 858 43240 13450 43352
rect 13618 43240 15384 43352
rect 858 43210 15384 43240
rect 858 43208 868 43210
rect 7108 43026 7240 43031
rect 7108 43020 7118 43026
rect 1036 42820 1046 43020
rect 1246 42914 7118 43020
rect 7230 43020 7240 43026
rect 7230 42914 7266 43020
rect 1246 42820 7266 42914
rect 12036 41478 12244 41483
rect 12036 41298 12046 41478
rect 12234 41298 12244 41478
rect 12036 41293 12244 41298
rect 6362 23314 6682 23319
rect 6362 23014 6372 23314
rect 6672 23014 6682 23314
rect 6362 23009 6682 23014
rect 106 22466 116 22974
rect 524 22882 554 22974
rect 1494 22882 1814 22887
rect 524 22582 1504 22882
rect 1804 22582 1814 22882
rect 524 22466 554 22582
rect 1494 22577 1814 22582
<< via3 >>
rect 14044 44738 14108 44818
rect 14596 44738 14660 44818
rect 15148 44738 15212 44818
rect 14950 43900 14952 43980
rect 14952 43900 15012 43980
rect 15012 43900 15014 43980
rect 9171 43724 9277 43729
rect 9171 43628 9176 43724
rect 9176 43628 9272 43724
rect 9272 43628 9277 43724
rect 9171 43623 9277 43628
rect 658 43208 858 43408
rect 1046 42820 1246 43020
rect 12046 41298 12234 41478
rect 6372 23014 6672 23314
rect 116 22466 524 22974
<< metal4 >>
rect 3006 45012 3066 45152
rect 3558 45012 3618 45152
rect 4110 45012 4170 45152
rect 4662 45012 4722 45152
rect 5214 45012 5274 45152
rect 5766 45012 5826 45152
rect 6318 45012 6378 45152
rect 6870 45012 6930 45152
rect 7422 45012 7482 45152
rect 7974 45012 8034 45152
rect 8526 45012 8586 45152
rect 9078 45012 9138 45152
rect 9630 45012 9690 45152
rect 10182 45012 10242 45152
rect 10734 45012 10794 45152
rect 11286 45012 11346 45152
rect 11838 45012 11898 45152
rect 12390 45012 12450 45152
rect 12942 45012 13002 45152
rect 13494 45012 13554 45152
rect 3006 44952 13554 45012
rect 8888 44610 8948 44952
rect 14046 44819 14106 45152
rect 14598 44819 14658 45152
rect 15150 44819 15210 45152
rect 14043 44818 14109 44819
rect 14043 44738 14044 44818
rect 14108 44738 14109 44818
rect 14043 44737 14109 44738
rect 14595 44818 14661 44819
rect 14595 44738 14596 44818
rect 14660 44738 14661 44818
rect 14595 44737 14661 44738
rect 15147 44818 15213 44819
rect 15147 44738 15148 44818
rect 15212 44738 15213 44818
rect 15147 44737 15213 44738
rect 200 44410 9170 44610
rect 15702 44422 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 200 22975 500 44410
rect 600 43408 900 44152
rect 600 43208 658 43408
rect 858 43208 900 43408
rect 115 22974 538 22975
rect 115 22466 116 22974
rect 524 22466 538 22974
rect 115 22465 538 22466
rect 200 1000 500 22465
rect 600 1000 900 43208
rect 1000 43020 1300 44152
rect 8970 43730 9170 44410
rect 14954 44362 15762 44422
rect 14954 44000 15014 44362
rect 14932 43980 15032 44000
rect 14932 43900 14950 43980
rect 15014 43900 15032 43980
rect 14932 43880 15032 43900
rect 8970 43729 9278 43730
rect 8970 43628 9171 43729
rect 9170 43623 9171 43628
rect 9277 43623 9278 43729
rect 9170 43622 9278 43623
rect 14954 43566 15014 43880
rect 1000 42820 1046 43020
rect 1246 42820 1300 43020
rect 1000 23314 1300 42820
rect 12045 41478 12235 41479
rect 12045 41298 12046 41478
rect 12234 41370 12235 41478
rect 28702 41370 28762 41374
rect 12234 41310 28762 41370
rect 12234 41298 12235 41310
rect 12045 41297 12235 41298
rect 6371 23314 6673 23315
rect 1000 23014 6372 23314
rect 6672 23014 6673 23314
rect 1000 1000 1300 23014
rect 6371 23013 6673 23014
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27234 198 27414 234
rect 28702 198 28762 41310
rect 27234 138 28762 198
rect 27234 0 27414 138
use big_skull  big_skull_0
timestamp 1735637413
transform 1 0 9298 0 1 31892
box 884 -15028 10166 -1768
use freq_divider  freq_divider_0
timestamp 1735637413
transform -1 0 18944 0 1 43628
box 3864 0 9552 640
use ring  ring_0
timestamp 1735637413
transform 1 0 14888 0 1 22922
box -12872 -12872 12872 12872
use skullfet_inverter_5v  skullfet_3v3_buffer
timestamp 1735637413
transform 0 1 7310 -1 0 43580
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_level_shifter
timestamp 1735637413
transform 0 -1 13802 -1 0 43580
box 454 132 2110 3088
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 43 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 44 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 45 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 46 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 47 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 48 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 49 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 50 nsew signal bidirectional
flabel metal4 1000 1000 1300 44152 1 FreeSans 2 0 0 0 VAPWR
port 51 nsew power bidirectional
flabel metal4 600 1000 900 44152 1 FreeSans 2 0 0 0 VDPWR
port 52 nsew power bidirectional
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VGND
port 53 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
