magic
tech sky130A
magscale 1 2
timestamp 1735290363
<< nwell >>
rect 676 132 1832 1400
<< pwell >>
rect 676 1944 1832 3088
<< mvnmos >>
rect 810 2619 1710 2719
<< mvpmos >>
rect 810 561 1710 661
<< mvndiff >>
rect 1050 2954 1530 3014
rect 990 2894 1530 2954
rect 870 2876 1650 2894
rect 870 2810 888 2876
rect 932 2810 1650 2876
rect 870 2774 1650 2810
rect 810 2719 1710 2774
rect 810 2566 1710 2619
rect 810 2500 822 2566
rect 866 2534 1710 2566
rect 866 2500 990 2534
rect 810 2474 990 2500
rect 810 2414 930 2474
rect 870 2354 930 2414
rect 1170 2354 1350 2534
rect 1530 2474 1710 2534
rect 1590 2414 1710 2474
rect 1590 2354 1650 2414
rect 870 2294 990 2354
rect 1110 2294 1410 2354
rect 1530 2294 1650 2354
rect 870 2234 1230 2294
rect 1290 2234 1590 2294
rect 990 2174 1170 2234
rect 1350 2174 1590 2234
rect 1050 2054 1470 2174
rect 1050 1994 1110 2054
rect 1170 1994 1230 2054
rect 1290 1994 1350 2054
rect 1410 1994 1470 2054
<< mvpdiff >>
rect 1050 1214 1110 1274
rect 1170 1214 1230 1274
rect 1290 1214 1350 1274
rect 1410 1214 1470 1274
rect 1050 1094 1470 1214
rect 990 1034 1170 1094
rect 1350 1034 1590 1094
rect 870 974 1230 1034
rect 1290 974 1590 1034
rect 870 914 990 974
rect 1110 914 1410 974
rect 1530 914 1650 974
rect 870 854 930 914
rect 810 794 930 854
rect 810 766 990 794
rect 810 700 822 766
rect 888 734 990 766
rect 1170 734 1350 914
rect 1590 854 1650 914
rect 1590 794 1710 854
rect 1530 734 1710 794
rect 888 700 1710 734
rect 810 661 1710 700
rect 810 494 1710 561
rect 870 454 1650 494
rect 870 388 888 454
rect 932 388 1650 454
rect 870 374 1650 388
rect 990 314 1530 374
rect 1050 254 1530 314
<< mvndiffc >>
rect 888 2810 932 2876
rect 822 2500 866 2566
<< mvpdiffc >>
rect 822 700 888 766
rect 888 388 932 454
<< mvpsubdiff >>
rect 732 3054 910 3066
rect 732 2972 766 3054
rect 876 2972 910 3054
<< mvnsubdiff >>
rect 744 300 900 310
rect 744 222 776 300
rect 866 222 900 300
rect 744 210 900 222
<< mvpsubdiffcont >>
rect 766 2972 876 3054
<< mvnsubdiffcont >>
rect 776 222 866 300
<< poly >>
rect 554 2619 810 2719
rect 1710 2619 2000 2719
rect 1888 2166 2000 2619
rect 1888 2054 1910 2166
rect 1976 2054 2000 2166
rect 1888 1188 2000 2054
rect 1888 1076 1910 1188
rect 1976 1076 2000 1188
rect 1888 661 2000 1076
rect 554 561 810 661
rect 1710 561 2000 661
<< polycont >>
rect 1910 2054 1976 2166
rect 1910 1076 1976 1188
<< locali >>
rect 732 3054 910 3066
rect 732 2972 766 3054
rect 876 2972 910 3054
rect 732 2900 910 2972
rect 688 2876 954 2900
rect 688 2822 710 2876
rect 766 2822 888 2876
rect 688 2810 888 2822
rect 932 2810 954 2876
rect 688 2788 954 2810
rect 554 2566 888 2588
rect 554 2500 822 2566
rect 866 2500 888 2566
rect 554 2476 888 2500
rect 554 1732 666 2476
rect 554 1576 566 1732
rect 654 1576 666 1732
rect 554 788 666 1576
rect 1888 2166 2000 2210
rect 1888 2054 1910 2166
rect 1976 2054 2000 2166
rect 1888 1732 2000 2054
rect 1888 1576 1900 1732
rect 1988 1576 2000 1732
rect 1888 1188 2000 1576
rect 1888 1076 1910 1188
rect 1976 1076 2000 1188
rect 1888 1010 2000 1076
rect 554 766 910 788
rect 554 700 822 766
rect 888 700 910 766
rect 554 676 910 700
rect 754 454 954 476
rect 754 432 888 454
rect 754 388 766 432
rect 822 388 888 432
rect 932 388 954 454
rect 754 366 954 388
rect 744 300 900 366
rect 744 222 776 300
rect 866 222 900 300
rect 744 210 900 222
<< viali >>
rect 710 2822 766 2876
rect 566 1576 654 1732
rect 1900 1576 1988 1732
rect 766 388 822 432
<< metal1 >>
rect 1050 2954 1530 3014
rect 554 2900 644 2922
rect 554 2822 566 2900
rect 632 2876 776 2900
rect 990 2894 1530 2954
rect 632 2822 710 2876
rect 766 2822 776 2876
rect 554 2800 776 2822
rect 870 2774 1650 2894
rect 810 2534 1710 2774
rect 810 2474 990 2534
rect 810 2414 930 2474
rect 870 2354 930 2414
rect 1170 2354 1350 2534
rect 1530 2474 1710 2534
rect 1590 2414 1710 2474
rect 1590 2354 1650 2414
rect 870 2294 990 2354
rect 1110 2294 1410 2354
rect 1530 2294 1650 2354
rect 870 2234 1230 2294
rect 1290 2234 1590 2294
rect 990 2174 1170 2234
rect 1350 2174 1590 2234
rect 1050 2054 1470 2174
rect 690 1994 870 2054
rect 1050 1994 1110 2054
rect 1170 1994 1230 2054
rect 1290 1994 1350 2054
rect 1410 1994 1470 2054
rect 1650 1994 1830 2054
rect 630 1874 930 1994
rect 1590 1874 1890 1994
rect 690 1814 1050 1874
rect 1470 1814 1830 1874
rect 870 1754 1110 1814
rect 1410 1754 1650 1814
rect 454 1732 666 1754
rect 454 1576 566 1732
rect 654 1576 666 1732
rect 990 1694 1230 1754
rect 1290 1694 1530 1754
rect 1888 1732 2110 1754
rect 454 1554 666 1576
rect 1110 1574 1410 1694
rect 1888 1576 1900 1732
rect 1988 1576 2110 1732
rect 990 1514 1230 1574
rect 1290 1514 1530 1574
rect 1888 1554 2110 1576
rect 690 1454 1110 1514
rect 1410 1454 1890 1514
rect 630 1394 990 1454
rect 1530 1394 1890 1454
rect 630 1334 870 1394
rect 1650 1334 1890 1394
rect 630 1274 810 1334
rect 1710 1274 1890 1334
rect 690 1214 750 1274
rect 1050 1214 1110 1274
rect 1170 1214 1230 1274
rect 1290 1214 1350 1274
rect 1410 1214 1470 1274
rect 1770 1214 1830 1274
rect 1050 1094 1470 1214
rect 990 1034 1170 1094
rect 1350 1034 1590 1094
rect 870 974 1230 1034
rect 1290 974 1590 1034
rect 870 914 990 974
rect 1110 914 1410 974
rect 1530 914 1650 974
rect 870 854 930 914
rect 810 794 930 854
rect 810 734 990 794
rect 1170 734 1350 914
rect 1590 854 1650 914
rect 1590 794 1710 854
rect 1530 734 1710 794
rect 810 494 1710 734
rect 554 432 832 454
rect 554 354 566 432
rect 654 388 766 432
rect 822 388 832 432
rect 654 366 832 388
rect 870 374 1650 494
rect 654 354 666 366
rect 554 332 666 354
rect 990 314 1530 374
rect 1050 254 1530 314
<< via1 >>
rect 566 2822 632 2900
rect 566 354 654 432
<< metal2 >>
rect 554 2900 644 3088
rect 1050 2954 1530 3014
rect 554 2822 566 2900
rect 632 2822 644 2900
rect 990 2894 1530 2954
rect 554 2800 644 2822
rect 870 2774 1650 2894
rect 810 2534 1710 2774
rect 810 2474 990 2534
rect 810 2414 930 2474
rect 870 2354 930 2414
rect 1170 2354 1350 2534
rect 1530 2474 1710 2534
rect 1590 2414 1710 2474
rect 1590 2354 1650 2414
rect 870 2294 990 2354
rect 1110 2294 1410 2354
rect 1530 2294 1650 2354
rect 870 2234 1230 2294
rect 1290 2234 1590 2294
rect 990 2174 1170 2234
rect 1350 2174 1590 2234
rect 1050 2054 1470 2174
rect 690 1994 870 2054
rect 1050 1994 1110 2054
rect 1170 1994 1230 2054
rect 1290 1994 1350 2054
rect 1410 1994 1470 2054
rect 1650 1994 1830 2054
rect 630 1874 930 1994
rect 1590 1874 1890 1994
rect 690 1814 1050 1874
rect 1470 1814 1830 1874
rect 870 1754 1110 1814
rect 1410 1754 1650 1814
rect 990 1694 1230 1754
rect 1290 1694 1530 1754
rect 1110 1574 1410 1694
rect 990 1514 1230 1574
rect 1290 1514 1530 1574
rect 690 1454 1110 1514
rect 1410 1454 1890 1514
rect 630 1394 990 1454
rect 1530 1394 1890 1454
rect 630 1334 870 1394
rect 1650 1334 1890 1394
rect 630 1274 810 1334
rect 1710 1274 1890 1334
rect 690 1214 750 1274
rect 1050 1214 1110 1274
rect 1170 1214 1230 1274
rect 1290 1214 1350 1274
rect 1410 1214 1470 1274
rect 1770 1214 1830 1274
rect 1050 1094 1470 1214
rect 990 1034 1170 1094
rect 1350 1034 1590 1094
rect 870 974 1230 1034
rect 1290 974 1590 1034
rect 870 914 990 974
rect 1110 914 1410 974
rect 1530 914 1650 974
rect 870 854 930 914
rect 810 794 930 854
rect 810 734 990 794
rect 1170 734 1350 914
rect 1590 854 1650 914
rect 1590 794 1710 854
rect 1530 734 1710 794
rect 810 494 1710 734
rect 554 432 666 454
rect 554 354 566 432
rect 654 354 666 432
rect 870 374 1650 494
rect 554 176 666 354
rect 990 314 1530 374
rect 1050 254 1530 314
<< obsm3 >>
rect 576 176 1954 3088
<< fillblock >>
rect 576 176 1954 3088
<< labels >>
flabel metal1 s 554 2800 644 2900 0 FreeSans 480 90 0 0 VGND
port 1 nsew ground bidirectional abutment
flabel metal1 s 554 366 666 454 0 FreeSans 480 90 0 0 VPWR
port 2 nsew power bidirectional abutment
flabel locali s 554 1566 666 1744 0 FreeSans 680 0 0 0 Y
port 3 s signal output
flabel locali s 1888 1566 2000 1744 0 FreeSans 680 0 0 0 A
port 4 e signal input
<< end >>
