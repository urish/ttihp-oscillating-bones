* NGSPICE file created from tt_um_oscillating_bones.ext - technology: ihp-sg13g2

.subckt tt_um_oscillating_bones ena clk rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] VGND VDPWR
X0 uo_out[1].t1 a_22205_61585# VGND.t33 VGND.t32 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X1 VDPWR.t44 a_16367_61578# freq_divider_0.sg13g2_dfrbp_2_0.D VDPWR.t0 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X2 VGND.t28 a_17996_61559# a_17075_61640# VGND.t27 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X3 VGND.t116 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_21132_61704# VGND.t115 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X4 a_16707_61717# a_16367_61578# VDPWR.t44 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X5 a_17910_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t19 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X6 a_20876_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t36 VDPWR.t0 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X7 ring_0/inverter_ring_0/skullfet_inverter_19.A ring_0/inverter_ring_0/skullfet_inverter_0.Y VDPWR.t39 VDPWR.t38 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X8 VGND.t16 a_22511_61578# a_22205_61585# VGND.t20 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X9 VGND.t114 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_18252_61704# VGND.t113 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X10 ring_0/inverter_ring_0/skullfet_inverter_6.A ring_0/inverter_ring_0/skullfet_inverter_7.A VDPWR.t18 VDPWR.t17 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X11 VGND.t47 ring_0/inverter_ring_0/skullfet_inverter_13.A ring_0/inverter_ring_0/skullfet_inverter_12.A VGND.t46 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X12 VDPWR.t16 a_20876_61559# a_19955_61640# VDPWR.t0 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X13 a_23109_61717# a_22851_61717# VGND.t49 VGND.t48 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X14 a_24054_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t15 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X15 VGND.t121 ring_0/inverter_ring_0/skullfet_inverter_17.A ring_0/inverter_ring_0/skullfet_inverter_16.A VGND.t120 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X16 VGND.t14 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_16801_61717# VGND.t13 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X17 a_20876_61559# a_19947_61366# a_20747_61559# VGND.t1 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X18 ring_0/inverter_ring_0/skullfet_inverter_12.A ring_0/inverter_ring_0/skullfet_inverter_13.A VDPWR.t33 VDPWR.t32 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X19 VDPWR.t13 a_22511_61578# freq_divider_0.sg13g2_dfrbp_2_2.D VDPWR.t0 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X20 a_23211_61366# a_23350_61250# VDPWR.t23 VDPWR.t0 sg13_lv_pmos ad=0.3864p pd=2.93u as=1.55707p ps=9.54u w=1.12u l=0.13u
X21 a_23211_61366# a_23350_61250# VGND.t55 VGND.t54 sg13_lv_nmos ad=0.2516p pd=2.16u as=2.07232p ps=13.14u w=0.74u l=0.13u
X22 VGND.t94 ring_0/inverter_ring_0/skullfet_inverter_9.A ring_0/inverter_ring_0/skullfet_inverter_8.A VGND.t93 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X23 ring_0/inverter_ring_0/skullfet_inverter_11.A ring_0/inverter_ring_0/skullfet_inverter_12.A VDPWR.t25 VDPWR.t24 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X24 VDPWR.t51 freq_divider_0.sg13g2_dfrbp_2_2.D a_24054_61326# VDPWR.t0 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X25 a_22851_61717# a_22511_61578# VDPWR.t13 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X26 a_23161_61402# a_22851_61717# VDPWR.t23 VDPWR.t0 sg13_lv_pmos ad=52.5f pd=0.67u as=1.55707p ps=9.54u w=0.42u l=0.13u
X27 VDPWR.t42 a_16367_61578# a_16061_61585# VDPWR.t0 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X28 a_17996_61559# a_17067_61366# a_17867_61559# VGND.t81 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X29 freq_divider_0.sg13g2_dfrbp_2_1.D a_19247_61578# VDPWR.t68 VDPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X30 VDPWR.t23 a_21777_61520# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t0 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3927p ps=2.99u w=1.155u l=0.13u
X31 a_22945_61717# a_22511_61578# a_22851_61717# VGND.t19 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X32 VGND.t111 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_24396_61704# VGND.t110 sg13_lv_nmos ad=0.1701p pd=1.65u as=38.85f ps=0.605u w=0.42u l=0.13u
X33 VDPWR.t11 a_22511_61578# a_22205_61585# VDPWR.t0 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X34 ring_0/inverter_ring_0/skullfet_inverter_3.A ring_0/inverter_ring_0/skullfet_inverter_4.A VDPWR.t60 VDPWR.t59 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X35 a_24396_61704# a_23219_61640# a_24011_61559# VGND.t68 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X36 a_21856_61617# a_21980_61316# VDPWR.t23 VDPWR.t0 sg13_lv_pmos ad=0.2442p pd=2.06u as=1.55707p ps=9.54u w=0.66u l=0.13u
X37 uo_out[2].t1 a_18941_61585# VGND.t43 VGND.t42 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X38 ring_0/inverter_ring_0/skullfet_inverter_17.A ring_0/inverter_ring_0/skullfet_inverter_18.A VDPWR.t41 VDPWR.t40 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X39 VGND.t70 ring_0/inverter_ring_0/skullfet_inverter_14.A ring_0/inverter_ring_0/skullfet_inverter_13.A VGND.t69 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X40 uo_out[2].t0 a_18941_61585# VDPWR.t31 VDPWR.t0 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X41 VGND.t37 ring_0/inverter_ring_0/skullfet_inverter_2.A ring_0/inverter_ring_0/skullfet_inverter_1.A VGND.t36 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X42 a_19247_61578# a_19947_61366# a_19897_61402# VDPWR.t0 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X43 ring_0/inverter_ring_0/skullfet_inverter_4.A ring_0/inverter_ring_0/skullfet_inverter_5.A VDPWR.t73 VDPWR.t72 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X44 VGND.t12 ring_0/inverter_ring_0/skullfet_inverter_11.A ring_0/inverter_ring_0/skullfet_inverter_10.A VGND.t11 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X45 VDPWR.t30 a_18941_61585# uo_out[2].t0 VDPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X46 VGND.t5 ring_0/inverter_ring_0/skullfet_inverter_0.A ring_0/inverter_ring_0/skullfet_inverter_0.Y VGND.t4 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X47 a_20876_61559# a_19947_61366# a_20790_61326# VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X48 a_18106_61326# a_17206_61250# a_17996_61559# VDPWR.t0 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X49 VGND.t39 ring_0/inverter_ring_0/skullfet_inverter_3.A ring_0/inverter_ring_0/skullfet_inverter_2.A VGND.t38 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X50 VGND.t118 ring_0/inverter_ring_0/skullfet_inverter_16.A uo_out[0].t1 VGND.t117 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X51 ring_0/inverter_ring_0/skullfet_inverter_18.A ring_0/inverter_ring_0/skullfet_inverter_19.A VDPWR.t53 VDPWR.t52 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X52 a_19947_61366# a_20086_61250# VDPWR.t23 VDPWR.t0 sg13_lv_pmos ad=0.3864p pd=2.93u as=1.55707p ps=9.54u w=1.12u l=0.13u
X53 ring_0/inverter_ring_0/skullfet_inverter_9.A ring_0/inverter_ring_0/skullfet_inverter_10.A VDPWR.t58 VDPWR.t57 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X54 VGND.t18 a_22511_61578# freq_divider_0.sg13g2_dfrbp_2_2.D VGND.t17 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X55 VGND.t90 uo_out[0].t2 ring_0/inverter_ring_0/skullfet_inverter_14.A VGND.t89 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X56 VGND.t31 a_22205_61585# uo_out[1].t1 VGND.t30 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X57 a_19681_61717# a_19247_61578# a_19587_61717# VGND.t100 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X58 a_17996_61559# a_17067_61366# a_17910_61326# VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X59 a_19955_61640# a_20086_61250# a_19247_61578# VDPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X60 a_20986_61326# a_20086_61250# a_20876_61559# VDPWR.t0 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X61 VDPWR.t10 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_16707_61717# VDPWR.t0 sg13_lv_pmos ad=1.4373p pd=8.805u as=79.8f ps=0.8u w=0.42u l=0.13u
X62 a_24140_61559# a_23211_61366# a_24054_61326# VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.1428p ps=1.52u w=0.42u l=0.13u
X63 a_17067_61366# a_17206_61250# VDPWR.t10 VDPWR.t0 sg13_lv_pmos ad=0.3864p pd=2.93u as=1.55707p ps=9.54u w=1.12u l=0.13u
X64 VDPWR.t23 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_22851_61717# VDPWR.t0 sg13_lv_pmos ad=1.4373p pd=8.805u as=79.8f ps=0.8u w=0.42u l=0.13u
X65 a_17067_61366# a_17206_61250# VGND.t79 VGND.t78 sg13_lv_nmos ad=0.2516p pd=2.16u as=2.07232p ps=13.14u w=0.74u l=0.13u
X66 VDPWR.t35 freq_divider_0.sg13g2_dfrbp_2_0.D a_17910_61326# VDPWR.t0 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X67 freq_divider_0.sg13g2_dfrbp_2_1.D a_19247_61578# VGND.t96 VGND.t99 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X68 a_21132_61704# a_19955_61640# a_20747_61559# VGND.t51 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X69 a_17910_61326# a_17206_61250# a_17996_61559# VGND.t123 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X70 a_19845_61717# a_20086_61250# a_19247_61578# VGND.t88 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X71 a_16965_61717# a_16707_61717# VGND.t14 VGND.t13 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X72 a_19897_61402# a_19587_61717# VDPWR.t10 VDPWR.t0 sg13_lv_pmos ad=52.5f pd=0.67u as=1.55707p ps=9.54u w=0.42u l=0.13u
X73 a_20790_61326# a_20086_61250# a_20876_61559# VGND.t87 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X74 a_18252_61704# a_17075_61640# a_17867_61559# VGND.t8 sg13_lv_nmos ad=38.85f pd=0.605u as=0.1596p ps=1.6u w=0.42u l=0.13u
X75 VGND.t98 a_19247_61578# freq_divider_0.sg13g2_dfrbp_2_1.D VGND.t97 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X76 VGND.t41 a_18941_61585# uo_out[2].t1 VGND.t40 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X77 a_24140_61559# a_23211_61366# a_24011_61559# VGND.t45 sg13_lv_nmos ad=81f pd=0.81u as=0.2163p ps=1.87u w=0.42u l=0.13u
X78 a_16965_61717# a_17206_61250# a_16367_61578# VGND.t122 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X79 VGND.t96 a_19247_61578# a_18941_61585# VGND.t95 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X80 a_17996_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t5 VDPWR.t0 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X81 VDPWR.t36 a_19955_61640# a_20986_61326# VDPWR.t0 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X82 a_20790_61326# freq_divider_0.sg13g2_dfrbp_2_1.D a_21529_61717# VGND.t29 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X83 VDPWR.t19 a_17996_61559# a_17075_61640# VDPWR.t0 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X84 VGND.t57 ring_0/inverter_ring_0/skullfet_inverter_0.Y ring_0/inverter_ring_0/skullfet_inverter_19.A VGND.t56 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X85 a_24140_61559# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t48 VDPWR.t0 sg13_lv_pmos ad=0.147p pd=1.54u as=0.1563p ps=1.22u w=0.42u l=0.13u
X86 ring_0/inverter_ring_0/skullfet_inverter_5.A ring_0/inverter_ring_0/skullfet_inverter_6.A VDPWR.t7 VDPWR.t6 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X87 VDPWR.t69 a_19247_61578# freq_divider_0.sg13g2_dfrbp_2_1.D VDPWR.t0 sg13_lv_pmos ad=0.2014p pd=1.53u as=0.2128p ps=1.5u w=1.12u l=0.13u
X88 VGND.t3 ring_0/inverter_ring_0/skullfet_inverter_8.A ring_0/inverter_ring_0/skullfet_inverter_7.A VGND.t2 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X89 VDPWR.t23 uo_out[1].t2 a_20086_61250# VDPWR.t0 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3808p ps=2.92u w=1.12u l=0.13u
X90 VDPWR.t15 a_24140_61559# a_23219_61640# VDPWR.t0 sg13_lv_pmos ad=0.36237p pd=2.605u as=0.34p ps=2.68u w=1u l=0.13u
X91 a_23219_61640# a_23350_61250# a_22511_61578# VDPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X92 VDPWR.t5 a_17075_61640# a_18106_61326# VDPWR.t0 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X93 a_19587_61717# a_19247_61578# VDPWR.t69 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.2014p ps=1.53u w=0.42u l=0.13u
X94 VGND.t67 ring_0/inverter_ring_0/skullfet_inverter_1.A ring_0/inverter_ring_0/skullfet_inverter_0.A VGND.t66 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X95 ring_0/inverter_ring_0/skullfet_inverter_10.A ring_0/inverter_ring_0/skullfet_inverter_11.A VDPWR.t9 VDPWR.t8 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X96 VDPWR.t22 a_22205_61585# uo_out[1].t0 VDPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X97 VDPWR.t10 uo_out[2].t2 a_17206_61250# VDPWR.t0 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3808p ps=2.92u w=1.12u l=0.13u
X98 VGND.t35 ring_0/inverter_ring_0/skullfet_inverter_12.A ring_0/inverter_ring_0/skullfet_inverter_11.A VGND.t34 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X99 a_23109_61717# a_23350_61250# a_22511_61578# VGND.t53 sg13_lv_nmos ad=0.1428p pd=1.52u as=0.12665p ps=1.145u w=0.42u l=0.13u
X100 ring_0/inverter_ring_0/skullfet_inverter_0.A ring_0/inverter_ring_0/skullfet_inverter_1.A VDPWR.t47 VDPWR.t46 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X101 ring_0/inverter_ring_0/skullfet_inverter_16.A ring_0/inverter_ring_0/skullfet_inverter_17.A VDPWR.t88 VDPWR.t87 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X102 a_21980_61316# a_21980_61316# VGND.t7 VGND.t92 sg13_lv_nmos ad=0.111p pd=1.34u as=2.07232p ps=13.14u w=0.3u l=0.13u
X103 VGND.t109 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_19681_61717# VGND.t108 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X104 ring_0/inverter_ring_0/skullfet_inverter_2.A ring_0/inverter_ring_0/skullfet_inverter_3.A VDPWR.t29 VDPWR.t28 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X105 uo_out[0].t0 ring_0/inverter_ring_0/skullfet_inverter_16.A VDPWR.t84 VDPWR.t83 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X106 a_21529_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t24 VGND.t107 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X107 VGND.t24 a_20876_61559# a_19955_61640# VGND.t23 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X108 uo_out[3].t1 a_16061_61585# VGND.t77 VGND.t76 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.2516p ps=2.16u w=0.74u l=0.13u
X109 VGND.t7 uo_out[1].t2 a_20086_61250# VGND.t6 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.2516p ps=2.16u w=0.74u l=0.13u
X110 VGND.t7 a_21856_61617# a_21777_61520# VGND.t101 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.27427p ps=2.28u w=0.795u l=0.13u
X111 a_16367_61578# a_17067_61366# a_17017_61402# VDPWR.t0 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X112 ring_0/inverter_ring_0/skullfet_inverter_14.A uo_out[0].t2 VDPWR.t63 VDPWR.t62 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X113 VGND.t85 ring_0/inverter_ring_0/skullfet_inverter_4.A ring_0/inverter_ring_0/skullfet_inverter_3.A VGND.t84 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X114 VDPWR.t48 a_23219_61640# a_24250_61326# VDPWR.t0 sg13_lv_pmos ad=0.1563p pd=1.22u as=54.6f ps=0.68u w=0.42u l=0.13u
X115 a_24250_61326# a_23350_61250# a_24140_61559# VDPWR.t0 sg13_lv_pmos ad=54.6f pd=0.68u as=79.8f ps=0.8u w=0.42u l=0.13u
X116 a_20790_61326# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VDPWR.t16 VDPWR.t0 sg13_lv_pmos ad=79.8f pd=0.8u as=0.36237p ps=2.605u w=0.42u l=0.13u
X117 a_24054_61326# freq_divider_0.sg13g2_dfrbp_2_2.D a_24793_61717# VGND.t71 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X118 a_22511_61578# a_23211_61366# a_23219_61640# VGND.t44 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X119 a_18649_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t28 VGND.t106 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X120 freq_divider_0.sg13g2_dfrbp_2_0.D a_16367_61578# VDPWR.t42 VDPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X121 VGND.t79 uo_out[2].t2 a_17206_61250# VGND.t78 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.2516p ps=2.16u w=0.74u l=0.13u
X122 VDPWR.t68 a_19247_61578# a_18941_61585# VDPWR.t0 sg13_lv_pmos ad=0.2083p pd=1.5u as=0.34p ps=2.68u w=1u l=0.13u
X123 VGND.t26 ring_0/inverter_ring_0/skullfet_inverter_7.A ring_0/inverter_ring_0/skullfet_inverter_6.A VGND.t25 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X124 a_24793_61717# freq_divider_0.sg13g2_dfrbp_2_0.RESET_B VGND.t22 VGND.t105 sg13_lv_nmos ad=60.89999f pd=0.71u as=0.1626p ps=1.415u w=0.42u l=0.13u
X125 a_17075_61640# a_17206_61250# a_16367_61578# VDPWR.t0 sg13_lv_pmos ad=0.34p pd=2.68u as=0.19115p ps=1.565u w=1u l=0.13u
X126 uo_out[3].t0 a_16061_61585# VDPWR.t55 VDPWR.t0 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X127 a_24054_61326# a_23350_61250# a_24140_61559# VGND.t52 sg13_lv_nmos ad=0.1296p pd=1.52u as=81f ps=0.81u w=0.42u l=0.13u
X128 VDPWR.t54 a_16061_61585# uo_out[3].t0 VDPWR.t0 sg13_lv_pmos ad=0.3808p pd=2.92u as=0.2156p ps=1.505u w=1.12u l=0.13u
X129 a_22511_61578# a_23211_61366# a_23161_61402# VDPWR.t0 sg13_lv_pmos ad=0.19115p pd=1.565u as=52.5f ps=0.67u w=0.42u l=0.13u
X130 ring_0/inverter_ring_0/skullfet_inverter_8.A ring_0/inverter_ring_0/skullfet_inverter_9.A VDPWR.t67 VDPWR.t66 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X131 uo_out[1].t0 a_22205_61585# VDPWR.t21 VDPWR.t0 sg13_lv_pmos ad=0.2156p pd=1.505u as=0.3808p ps=2.92u w=1.12u l=0.13u
X132 ring_0/inverter_ring_0/skullfet_inverter_7.A ring_0/inverter_ring_0/skullfet_inverter_8.A VDPWR.t2 VDPWR.t1 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X133 VGND.t83 ring_0/inverter_ring_0/skullfet_inverter_10.A ring_0/inverter_ring_0/skullfet_inverter_9.A VGND.t82 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X134 VGND.t22 a_24140_61559# a_23219_61640# VGND.t21 sg13_lv_nmos ad=0.1626p pd=1.415u as=0.2516p ps=2.16u w=0.74u l=0.13u
X135 VGND.t55 uo_out[0].t3 a_23350_61250# VGND.t54 sg13_lv_nmos ad=2.07232p pd=13.14u as=0.2516p ps=2.16u w=0.74u l=0.13u
X136 freq_divider_0.sg13g2_dfrbp_2_2.D a_22511_61578# VDPWR.t11 VDPWR.t0 sg13_lv_pmos ad=0.2128p pd=1.5u as=0.2083p ps=1.5u w=1.12u l=0.13u
X137 a_16801_61717# a_16367_61578# a_16707_61717# VGND.t65 sg13_lv_nmos ad=37.8f pd=0.6u as=0.1428p ps=1.52u w=0.42u l=0.13u
X138 a_19247_61578# a_19947_61366# a_19955_61640# VGND.t0 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X139 ring_0/inverter_ring_0/skullfet_inverter_1.A ring_0/inverter_ring_0/skullfet_inverter_2.A VDPWR.t27 VDPWR.t26 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X140 ring_0/inverter_ring_0/skullfet_inverter_13.A ring_0/inverter_ring_0/skullfet_inverter_14.A VDPWR.t50 VDPWR.t49 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X141 VDPWR.t10 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_19587_61717# VDPWR.t0 sg13_lv_pmos ad=1.4373p pd=8.805u as=79.8f ps=0.8u w=0.42u l=0.13u
X142 ring_0/inverter_ring_0/skullfet_inverter_0.Y ring_0/inverter_ring_0/skullfet_inverter_0.A VDPWR.t4 VDPWR.t3 sg13_lv_pmos ad=6.2694p pd=26.64u as=4.4307p ps=10.9u w=4.05u l=0.4u
X143 freq_divider_0.sg13g2_dfrbp_2_0.D a_16367_61578# VGND.t61 VGND.t64 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
X144 a_17910_61326# freq_divider_0.sg13g2_dfrbp_2_0.D a_18649_61717# VGND.t50 sg13_lv_nmos ad=0.1428p pd=1.52u as=60.89999f ps=0.71u w=0.42u l=0.13u
X145 a_16367_61578# a_17067_61366# a_17075_61640# VGND.t80 sg13_lv_nmos ad=0.12665p pd=1.145u as=0.3473p ps=2.71u w=0.74u l=0.13u
X146 VGND.t49 freq_divider_0.sg13g2_dfrbp_2_0.RESET_B a_22945_61717# VGND.t48 sg13_lv_nmos ad=79.8f pd=0.8u as=37.8f ps=0.6u w=0.42u l=0.13u
X147 a_17017_61402# a_16707_61717# VDPWR.t10 VDPWR.t0 sg13_lv_pmos ad=52.5f pd=0.67u as=1.55707p ps=9.54u w=0.42u l=0.13u
X148 VGND.t59 ring_0/inverter_ring_0/skullfet_inverter_18.A ring_0/inverter_ring_0/skullfet_inverter_17.A VGND.t58 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X149 VGND.t63 a_16367_61578# freq_divider_0.sg13g2_dfrbp_2_0.D VGND.t62 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X150 VGND.t10 ring_0/inverter_ring_0/skullfet_inverter_6.A ring_0/inverter_ring_0/skullfet_inverter_5.A VGND.t9 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X151 VGND.t75 a_16061_61585# uo_out[3].t1 VGND.t74 sg13_lv_nmos ad=0.2516p pd=2.16u as=0.1406p ps=1.12u w=0.74u l=0.13u
X152 a_19845_61717# a_19587_61717# VGND.t109 VGND.t108 sg13_lv_nmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X153 VGND.t103 ring_0/inverter_ring_0/skullfet_inverter_5.A ring_0/inverter_ring_0/skullfet_inverter_4.A VGND.t102 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X154 VGND.t61 a_16367_61578# a_16061_61585# VGND.t60 sg13_lv_nmos ad=0.1331p pd=1.12u as=0.2176p ps=1.96u w=0.64u l=0.13u
X155 VDPWR.t23 uo_out[0].t3 a_23350_61250# VDPWR.t0 sg13_lv_pmos ad=1.55707p pd=9.54u as=0.3808p ps=2.92u w=1.12u l=0.13u
X156 a_19947_61366# a_20086_61250# VGND.t7 VGND.t6 sg13_lv_nmos ad=0.2516p pd=2.16u as=2.07232p ps=13.14u w=0.74u l=0.13u
X157 VGND.t73 ring_0/inverter_ring_0/skullfet_inverter_19.A ring_0/inverter_ring_0/skullfet_inverter_18.A VGND.t72 sg13_lv_nmos ad=4.2687p pd=10.82u as=6.4314p ps=26.72u w=4.05u l=0.4u
X158 VDPWR.t20 freq_divider_0.sg13g2_dfrbp_2_1.D a_20790_61326# VDPWR.t0 sg13_lv_pmos ad=0.1428p pd=1.52u as=79.8f ps=0.8u w=0.42u l=0.13u
X159 freq_divider_0.sg13g2_dfrbp_2_2.D a_22511_61578# VGND.t16 VGND.t15 sg13_lv_nmos ad=0.1406p pd=1.12u as=0.1331p ps=1.12u w=0.74u l=0.13u
R0 VGND.n199 VGND.n59 36337.9
R1 VGND.n207 VGND.n111 26006.8
R2 VGND.n343 VGND.n111 20289.4
R3 VGND.t84 VGND.n157 19416.2
R4 VGND.n466 VGND.n465 17662.9
R5 VGND.n191 VGND.n70 15262.5
R6 VGND.n199 VGND.n111 12285.4
R7 VGND.n61 VGND.n59 12285.4
R8 VGND.n465 VGND.n464 12279.6
R9 VGND.n197 VGND.t9 12039.2
R10 VGND.t25 VGND.n63 10402.1
R11 VGND.n278 VGND.n271 10052.7
R12 VGND.n467 VGND.n466 10011.4
R13 VGND.n156 VGND.n155 9840.79
R14 VGND.n198 VGND.n61 9066.9
R15 VGND.n262 VGND.n197 7844.55
R16 VGND.n207 VGND.n201 7498.6
R17 VGND.n196 VGND.n195 7474.99
R18 VGND.n155 VGND.n152 7291.79
R19 VGND.n191 VGND.t102 7169.54
R20 VGND.n470 VGND.n65 6899.39
R21 VGND.n474 VGND.n60 6851.13
R22 VGND.n69 VGND.n65 6429.23
R23 VGND.n262 VGND.t38 6051.63
R24 VGND.n200 VGND.n199 6014.02
R25 VGND.n464 VGND.n463 5872.62
R26 VGND.n201 VGND.n200 5699.78
R27 VGND.n464 VGND.n69 5321.16
R28 VGND.n192 VGND.n191 5298.87
R29 VGND.n476 VGND.n475 4953.11
R30 VGND.n466 VGND.n69 4950.06
R31 VGND.n261 VGND.n260 4945.91
R32 VGND.n288 VGND.n152 3511.45
R33 VGND.n155 VGND.n154 3475.34
R34 VGND.n273 VGND.n268 3284.18
R35 VGND.n464 VGND.n71 3154.9
R36 VGND.n197 VGND.n196 3153.12
R37 VGND.n279 VGND.n278 2376.2
R38 VGND.n262 VGND.n154 2220.92
R39 VGND.n468 VGND.n467 2091.57
R40 VGND.n472 VGND.n63 1946.24
R41 VGND.n200 VGND.n198 1880.71
R42 VGND.n157 VGND.n70 1835.32
R43 VGND.n74 VGND.n71 1763.01
R44 VGND.n262 VGND.n198 1734.38
R45 VGND.n197 VGND.n63 1470.05
R46 VGND.n280 VGND.t4 1368.89
R47 VGND.t72 VGND.n273 1347.06
R48 VGND.n273 VGND.t56 1194.61
R49 VGND.t102 VGND.n190 1123.79
R50 VGND.n465 VGND.n70 1061.65
R51 VGND.n280 VGND.n268 977.779
R52 VGND.n60 VGND.t46 964.287
R53 VGND.n262 VGND.n156 905.553
R54 VGND.t46 VGND.n59 876.317
R55 VGND.n474 VGND.n61 837.723
R56 VGND.n272 VGND.n152 814.62
R57 VGND.n234 VGND.n231 744.615
R58 VGND.n484 VGND.n5 744.615
R59 VGND.n53 VGND.n52 744.615
R60 VGND.n206 VGND.t89 675.663
R61 VGND.n195 VGND.t38 656.004
R62 VGND.n463 VGND.t9 656.004
R63 VGND.n196 VGND.t84 615.229
R64 VGND.n156 VGND.n151 608.424
R65 VGND.n344 VGND.n59 575.212
R66 VGND.n196 VGND.n192 498.868
R67 VGND.n234 VGND.t48 480
R68 VGND.n484 VGND.t108 480
R69 VGND.n52 VGND.t13 480
R70 VGND.n469 VGND.t93 455.887
R71 VGND.n74 VGND.t25 427.755
R72 VGND.n262 VGND.n261 402.269
R73 VGND.n475 VGND.n474 395.865
R74 VGND.n262 VGND.n201 392.892
R75 VGND.t69 VGND.n343 372.399
R76 VGND.n279 VGND.n268 344.149
R77 VGND.t56 VGND.n271 335.173
R78 VGND.n68 VGND.t93 330.428
R79 VGND.n288 VGND.t120 318.406
R80 VGND.n343 VGND.n342 307.757
R81 VGND.n157 VGND.n154 278.079
R82 VGND.n230 VGND.t17 260.005
R83 VGND.n16 VGND.t97 260.005
R84 VGND.t62 VGND.n54 260.005
R85 VGND.t15 VGND.n228 234.738
R86 VGND.t99 VGND.n14 234.738
R87 VGND.n56 VGND.t64 234.738
R88 VGND.n241 VGND.t20 232.869
R89 VGND.n25 VGND.t95 232.869
R90 VGND.t60 VGND.n43 232.869
R91 VGND.t36 VGND.n151 231.615
R92 VGND.t101 VGND.n225 228.233
R93 VGND.n272 VGND.t66 227.947
R94 VGND.n198 VGND.n63 226.054
R95 VGND.n248 VGND.t23 200.339
R96 VGND.n31 VGND.t27 200.339
R97 VGND.n212 VGND.t21 200.339
R98 VGND.n246 VGND.t29 195.942
R99 VGND.n12 VGND.t50 194.969
R100 VGND.n473 VGND.n472 194.851
R101 VGND.n245 VGND.t30 185.124
R102 VGND.n29 VGND.t40 185.124
R103 VGND.t74 VGND.n41 185.124
R104 VGND.t32 VGND.n226 184.825
R105 VGND.t42 VGND.n12 184.825
R106 VGND.n260 VGND.t71 180.052
R107 VGND.n226 VGND.t92 172.145
R108 VGND.n476 VGND.t76 169.907
R109 VGND.n278 VGND.t58 164.255
R110 VGND.t51 VGND.t115 159.763
R111 VGND.t8 VGND.t113 159.763
R112 VGND.t68 VGND.t110 159.763
R113 VGND.t1 VGND.n221 156.929
R114 VGND.t81 VGND.n9 156.929
R115 VGND.t45 VGND.n209 156.929
R116 VGND.n252 VGND.t87 154.614
R117 VGND.n35 VGND.t123 154.614
R118 VGND.n215 VGND.t52 154.614
R119 VGND.n71 VGND.n65 151.276
R120 VGND.t107 VGND.n223 149.62
R121 VGND.t106 VGND.n11 149.62
R122 VGND.t105 VGND.n211 149.62
R123 VGND.t48 VGND.t44 138.463
R124 VGND.t108 VGND.t0 138.463
R125 VGND.t13 VGND.t80 138.463
R126 VGND.n261 VGND.t117 132.323
R127 VGND.n472 VGND.t2 128.216
R128 VGND.n475 VGND.n59 122.921
R129 VGND.t4 VGND.n279 113.026
R130 VGND.n231 VGND.t19 110.237
R131 VGND.t100 VGND.n5 110.237
R132 VGND.t65 VGND.n53 110.237
R133 VGND.n221 VGND.n5 106.212
R134 VGND.n53 VGND.n9 106.212
R135 VGND.n231 VGND.n209 106.212
R136 VGND.t87 VGND.n251 100.478
R137 VGND.t123 VGND.n34 100.478
R138 VGND.t52 VGND.n214 100.478
R139 VGND.n252 VGND.t1 99.7516
R140 VGND.n35 VGND.t81 99.7516
R141 VGND.n215 VGND.t45 99.7516
R142 VGND.n467 VGND.n68 95.8456
R143 VGND.t2 VGND.n471 95.5275
R144 VGND.n248 VGND.t107 93.8297
R145 VGND.n31 VGND.t106 93.8297
R146 VGND.n212 VGND.t105 93.8297
R147 VGND.t92 VGND.n225 86.222
R148 VGND.n288 VGND.n151 84.6642
R149 VGND.n471 VGND.n470 83.8532
R150 VGND.n251 VGND.t51 75.5501
R151 VGND.n34 VGND.t8 75.5501
R152 VGND.n214 VGND.t68 75.5501
R153 VGND.t54 VGND.t53 73.8467
R154 VGND.t6 VGND.t88 73.8467
R155 VGND.t78 VGND.t122 73.8467
R156 VGND.n245 VGND.t32 73.5423
R157 VGND.n29 VGND.t42 73.5423
R158 VGND.t76 VGND.n41 73.5423
R159 VGND.t30 VGND.n241 73.244
R160 VGND.t40 VGND.n25 73.244
R161 VGND.n43 VGND.t74 73.244
R162 VGND.n287 VGND.t66 72.396
R163 VGND.n342 VGND.t89 65.0575
R164 VGND.n344 VGND.t69 63.8663
R165 VGND.n474 VGND.t34 63.5677
R166 VGND.t29 VGND.n223 63.3986
R167 VGND.t50 VGND.n11 63.3986
R168 VGND.n211 VGND.t71 63.3986
R169 VGND.t21 VGND.n210 59.0031
R170 VGND.t23 VGND.n222 59.0031
R171 VGND.t27 VGND.n10 59.0031
R172 VGND.n472 VGND.t11 55.0827
R173 VGND.n263 VGND.t36 51.425
R174 VGND.n203 VGND.t120 51.1311
R175 VGND.t19 VGND.n230 48.4827
R176 VGND.n16 VGND.t100 48.4827
R177 VGND.n54 VGND.t65 48.4827
R178 VGND.t34 VGND.n473 47.9255
R179 VGND.n469 VGND.t82 47.7166
R180 VGND.n469 VGND.n66 44.7738
R181 VGND.n289 VGND.t58 44.7032
R182 VGND.t117 VGND.n207 42.4247
R183 VGND.n66 VGND.t11 41.6077
R184 VGND.n277 VGND.t72 38.7252
R185 VGND.t115 VGND.n222 38.7147
R186 VGND.t113 VGND.n10 38.7147
R187 VGND.t110 VGND.n210 38.7147
R188 VGND.n278 VGND.n272 36.6123
R189 VGND.t82 VGND.n468 36.1063
R190 VGND.n246 VGND.t101 31.1079
R191 VGND.t20 VGND.n228 28.3754
R192 VGND.t95 VGND.n14 28.3754
R193 VGND.n56 VGND.t60 28.3754
R194 VGND.n229 VGND.t15 27.8464
R195 VGND.n15 VGND.t99 27.8464
R196 VGND.t64 VGND.n55 27.8464
R197 VGND.t44 VGND.t54 24.6159
R198 VGND.t0 VGND.t6 24.6159
R199 VGND.t80 VGND.t78 24.6159
R200 VGND.n288 VGND.n287 22.6588
R201 VGND.n207 VGND.n206 22.6333
R202 VGND.n470 VGND.n469 18.8055
R203 VGND.n286 VGND.n285 18.1658
R204 VGND.n265 VGND.n264 18.1658
R205 VGND.n391 VGND.n390 18.1658
R206 VGND.n77 VGND.n64 18.1658
R207 VGND.n76 VGND.n75 18.1658
R208 VGND.n462 VGND.n461 18.1658
R209 VGND.n190 VGND.n189 18.1658
R210 VGND.n159 VGND.n158 18.1658
R211 VGND.n446 VGND.n445 18.1658
R212 VGND.n87 VGND.n67 18.1658
R213 VGND.n88 VGND.n62 18.1658
R214 VGND.n205 VGND.n204 18.1658
R215 VGND.n202 VGND.n140 18.1658
R216 VGND.n291 VGND.n290 18.1658
R217 VGND.n276 VGND.n275 18.1658
R218 VGND.n270 VGND.n269 18.1658
R219 VGND.n341 VGND.n340 18.1658
R220 VGND.n346 VGND.n345 18.1658
R221 VGND.n372 VGND.n371 18.1658
R222 VGND.n194 VGND.n193 18.1658
R223 VGND.n282 VGND.n281 18.1658
R224 VGND.t7 VGND.n252 18.0261
R225 VGND.t79 VGND.n35 18.0261
R226 VGND.t55 VGND.n215 18.0261
R227 VGND.t17 VGND.n229 17.5282
R228 VGND.t97 VGND.n15 17.5282
R229 VGND.n55 VGND.t62 17.5282
R230 VGND.n213 VGND.t22 17.2928
R231 VGND.n36 VGND.t114 17.2395
R232 VGND.n253 VGND.t116 17.2395
R233 VGND.n216 VGND.t111 17.2395
R234 VGND.n47 VGND.t63 17.2297
R235 VGND.n21 VGND.t98 17.2297
R236 VGND.n237 VGND.t18 17.2297
R237 VGND.n40 VGND.t14 17.2268
R238 VGND.n32 VGND.t28 17.2268
R239 VGND.n19 VGND.t109 17.2268
R240 VGND.n249 VGND.t24 17.2268
R241 VGND.n220 VGND.t49 17.2268
R242 VGND.n402 VGND.t61 17.212
R243 VGND.n23 VGND.t96 17.212
R244 VGND.n239 VGND.t16 17.212
R245 VGND.n57 VGND.t77 17.2025
R246 VGND.n27 VGND.t43 17.2025
R247 VGND.n243 VGND.t33 17.2025
R248 VGND.n286 VGND.t67 17.0362
R249 VGND.n264 VGND.t37 17.0362
R250 VGND.n390 VGND.t12 17.0362
R251 VGND.n64 VGND.t3 17.0362
R252 VGND.n75 VGND.t26 17.0362
R253 VGND.n462 VGND.t10 17.0362
R254 VGND.n190 VGND.t103 17.0362
R255 VGND.n158 VGND.t85 17.0362
R256 VGND.n445 VGND.t94 17.0362
R257 VGND.n67 VGND.t83 17.0362
R258 VGND.n62 VGND.t35 17.0362
R259 VGND.n205 VGND.t118 17.0362
R260 VGND.n202 VGND.t121 17.0362
R261 VGND.n290 VGND.t59 17.0362
R262 VGND.n276 VGND.t73 17.0362
R263 VGND.n270 VGND.t57 17.0362
R264 VGND.n341 VGND.t90 17.0362
R265 VGND.n345 VGND.t70 17.0362
R266 VGND.n371 VGND.t47 17.0362
R267 VGND.n194 VGND.t39 17.0362
R268 VGND.n281 VGND.t5 17.0362
R269 VGND.n260 VGND.t55 17.0005
R270 VGND.t55 VGND.n211 17.0005
R271 VGND.t55 VGND.n212 17.0005
R272 VGND.n255 VGND.t7 17.0005
R273 VGND.t7 VGND.n228 17.0005
R274 VGND.t7 VGND.n245 17.0005
R275 VGND.t7 VGND.n227 17.0005
R276 VGND.t7 VGND.n225 17.0005
R277 VGND.t7 VGND.n223 17.0005
R278 VGND.t7 VGND.n248 17.0005
R279 VGND.n486 VGND.n1 17.0005
R280 VGND.n487 VGND.n486 17.0005
R281 VGND.t79 VGND.n18 17.0005
R282 VGND.t79 VGND.n14 17.0005
R283 VGND.t79 VGND.n29 17.0005
R284 VGND.t79 VGND.n13 17.0005
R285 VGND.t79 VGND.n11 17.0005
R286 VGND.t79 VGND.n31 17.0005
R287 VGND.n478 VGND.n477 17.0005
R288 VGND.n477 VGND.n56 17.0005
R289 VGND.n477 VGND.n41 17.0005
R290 VGND.n477 VGND.n58 17.0005
R291 VGND.n477 VGND.n476 17.0005
R292 VGND.n281 VGND.n280 16.9935
R293 VGND.n263 VGND.n262 16.2915
R294 VGND.n262 VGND.n203 16.2014
R295 VGND.n468 VGND.n67 15.6652
R296 VGND.n277 VGND.n276 15.5838
R297 VGND.n390 VGND.n66 15.4962
R298 VGND.n290 VGND.n289 15.4044
R299 VGND.n473 VGND.n62 15.3111
R300 VGND.n203 VGND.n202 15.2207
R301 VGND.n264 VGND.n263 15.2126
R302 VGND.n345 VGND.n344 14.8829
R303 VGND.n206 VGND.n205 14.853
R304 VGND.n342 VGND.n341 14.853
R305 VGND.n287 VGND.n286 14.6742
R306 VGND.n289 VGND.n288 14.2225
R307 VGND.n471 VGND.n64 14.1685
R308 VGND.n278 VGND.n277 12.3693
R309 VGND.n489 VGND.n488 11.5981
R310 VGND.n404 VGND.n403 11.5903
R311 VGND.n445 VGND.n68 11.5621
R312 VGND.n271 VGND.n270 11.5336
R313 VGND.n75 VGND.n74 11.0666
R314 VGND.n463 VGND.n462 10.3577
R315 VGND.n195 VGND.n194 10.3577
R316 VGND.n371 VGND.n60 9.85117
R317 VGND.n192 VGND.n158 9.69267
R318 VGND.n433 VGND.n428 9.0005
R319 VGND.n428 VGND.n421 9.0005
R320 VGND.n433 VGND.n432 9.0005
R321 VGND.n432 VGND.n421 9.0005
R322 VGND.n433 VGND.n427 9.0005
R323 VGND.n434 VGND.n423 9.0005
R324 VGND.n434 VGND.n421 9.0005
R325 VGND.n434 VGND.n433 9.0005
R326 VGND.n439 VGND.n436 9.0005
R327 VGND.n436 VGND.n419 9.0005
R328 VGND.n439 VGND.n438 9.0005
R329 VGND.n438 VGND.n419 9.0005
R330 VGND.n439 VGND.n435 9.0005
R331 VGND.n441 VGND.n440 9.0005
R332 VGND.n440 VGND.n419 9.0005
R333 VGND.n440 VGND.n439 9.0005
R334 VGND.n440 uio_oe[7] 8.8478
R335 VGND.n44 VGND.t75 8.74885
R336 VGND.n26 VGND.t41 8.74885
R337 VGND.n242 VGND.t31 8.74885
R338 VGND.n234 VGND.n232 8.501
R339 VGND.n234 VGND.n233 8.501
R340 VGND.n485 VGND.n484 8.501
R341 VGND.n484 VGND.n6 8.501
R342 VGND.n52 VGND.n50 8.501
R343 VGND.n52 VGND.n51 8.501
R344 VGND.n258 VGND.n217 8.47111
R345 VGND.n257 VGND.n218 8.47111
R346 VGND.n256 VGND.n219 8.47111
R347 VGND.t7 VGND.n238 8.47111
R348 VGND.t7 VGND.n240 8.47111
R349 VGND.t7 VGND.n244 8.47111
R350 VGND.t7 VGND.n250 8.47111
R351 VGND.n4 VGND.n2 8.47111
R352 VGND.n17 VGND.n7 8.47111
R353 VGND.t79 VGND.n22 8.47111
R354 VGND.t79 VGND.n24 8.47111
R355 VGND.t79 VGND.n28 8.47111
R356 VGND.t79 VGND.n33 8.47111
R357 VGND.n481 VGND.n37 8.47111
R358 VGND.n480 VGND.n38 8.47111
R359 VGND.n479 VGND.n39 8.47111
R360 VGND.n477 VGND.n46 8.47111
R361 VGND.n477 VGND.n45 8.47111
R362 VGND.n477 VGND.n42 8.47111
R363 VGND.n266 VGND.n153 8.0799
R364 VGND.n458 VGND.n457 7.52168
R365 VGND.n458 VGND.n76 7.47272
R366 VGND.n274 VGND.n150 6.68645
R367 VGND.n461 VGND.n460 6.53659
R368 VGND.n160 VGND.n159 6.32858
R369 VGND.n392 VGND.n389 6.30123
R370 VGND.n189 VGND.n188 6.07977
R371 VGND.n193 VGND.n153 6.05718
R372 VGND.n266 VGND.n265 5.9638
R373 VGND.n235 VGND.n234 5.66778
R374 VGND.n484 VGND.n483 5.66778
R375 VGND.n52 VGND.n49 5.66778
R376 VGND.n234 VGND.n208 5.66767
R377 VGND.n484 VGND.n3 5.66767
R378 VGND.n52 VGND.n8 5.66767
R379 VGND.t7 VGND.n236 5.61485
R380 VGND.t7 VGND.n247 5.61485
R381 VGND.t79 VGND.n20 5.61485
R382 VGND.t79 VGND.n30 5.61485
R383 VGND.n477 VGND.n48 5.61485
R384 VGND.n284 VGND.n266 5.49409
R385 VGND.n427 VGND 5.4103
R386 VGND.n285 VGND.n284 4.52382
R387 VGND.n431 VGND.n430 4.49573
R388 VGND.n430 VGND.n422 4.49573
R389 VGND.n437 VGND.n394 4.49573
R390 VGND.n420 VGND.n394 4.49573
R391 VGND.n429 VGND.n423 4.49573
R392 VGND.n441 VGND.n397 4.49573
R393 VGND.n427 VGND.n426 4.4949
R394 VGND.n435 VGND.n396 4.4949
R395 VGND.n283 VGND.n282 4.09378
R396 VGND.n269 VGND.n267 3.42765
R397 VGND.t55 VGND.n213 3.38768
R398 VGND.t7 VGND.n224 3.34182
R399 VGND.n275 VGND.n274 3.27628
R400 VGND.n292 VGND.n291 2.85446
R401 VGND.n320 VGND.n125 2.31911
R402 VGND.n125 VGND 2.31911
R403 VGND.n78 VGND.n77 2.27849
R404 VGND.n443 VGND.n394 2.2505
R405 VGND.n442 VGND.n441 2.2505
R406 VGND.n430 VGND.n86 2.2505
R407 VGND.n424 VGND.n423 2.2505
R408 VGND.t55 VGND.n259 1.97699
R409 VGND.t7 VGND.n254 1.97699
R410 VGND.t79 VGND.n482 1.97699
R411 VGND.n447 VGND.n446 1.81263
R412 VGND.n306 VGND.n140 1.72671
R413 VGND.n340 VGND.n339 1.47805
R414 VGND.n339 VGND.n338 1.4745
R415 VGND.n435 VGND.n434 1.40696
R416 VGND.n393 VGND 1.31963
R417 VGND.t7 VGND.n251 1.21402
R418 VGND.t79 VGND.n34 1.21402
R419 VGND.t55 VGND.n214 1.21402
R420 VGND.n274 VGND.n267 1.18201
R421 VGND.n442 VGND.n395 1.1463
R422 VGND.n425 VGND.n424 1.1463
R423 VGND.n392 VGND.n391 1.13055
R424 VGND.t55 VGND.n209 1.04263
R425 VGND.t7 VGND.n241 1.04263
R426 VGND.t7 VGND.n226 1.04263
R427 VGND.t7 VGND.n221 1.04263
R428 VGND.t79 VGND.n25 1.04263
R429 VGND.t79 VGND.n12 1.04263
R430 VGND.t79 VGND.n9 1.04263
R431 VGND.n477 VGND.n43 1.04263
R432 VGND.t7 VGND.n230 1.02715
R433 VGND.t7 VGND.n229 1.02715
R434 VGND.t79 VGND.n16 1.02715
R435 VGND.t79 VGND.n15 1.02715
R436 VGND.n477 VGND.n54 1.02715
R437 VGND.n477 VGND.n55 1.02715
R438 VGND.n322 VGND.n125 0.936079
R439 VGND.n89 VGND.n88 0.882121
R440 VGND.n204 VGND.n125 0.851167
R441 VGND.n347 VGND.n346 0.8068
R442 VGND.n373 VGND.n372 0.803036
R443 VGND.n393 VGND.n392 0.620893
R444 VGND.n377 VGND.n376 0.598489
R445 VGND.n259 VGND.n258 0.585769
R446 VGND.n482 VGND.n481 0.585769
R447 VGND.n254 VGND.n1 0.52548
R448 VGND.n444 VGND.n443 0.521717
R449 VGND.n459 VGND.n458 0.518224
R450 VGND.n259 VGND.n216 0.477006
R451 VGND.n254 VGND.n253 0.477006
R452 VGND.n482 VGND.n36 0.477006
R453 VGND.n339 VGND.n112 0.473781
R454 VGND.n160 VGND.n153 0.464095
R455 VGND.n449 VGND.n86 0.45348
R456 VGND.n335 VGND.n112 0.434656
R457 VGND.n305 VGND.n141 0.423272
R458 VGND.n284 VGND.n283 0.364261
R459 VGND.n378 VGND.n377 0.352948
R460 VGND.n335 VGND.n334 0.347746
R461 VGND.n161 VGND.n160 0.328048
R462 VGND.n398 uo_out[5] 0.32522
R463 VGND.n399 uo_out[6] 0.32522
R464 VGND.n400 uo_out[7] 0.32522
R465 VGND.n401 uio_out[0] 0.32522
R466 VGND.n406 uio_out[2] 0.32522
R467 VGND.n407 uio_out[3] 0.32522
R468 VGND.n408 uio_out[4] 0.32522
R469 VGND.n409 uio_out[5] 0.32522
R470 VGND.n410 uio_out[6] 0.32522
R471 VGND.n411 uio_out[7] 0.32522
R472 VGND.n412 uio_oe[0] 0.32522
R473 VGND.n413 uio_oe[1] 0.32522
R474 VGND.n414 uio_oe[2] 0.32522
R475 VGND.n415 uio_oe[3] 0.32522
R476 VGND.n416 uio_oe[4] 0.32522
R477 VGND.n417 uio_oe[5] 0.32522
R478 VGND.n418 uio_oe[6] 0.32522
R479 VGND.n334 VGND.n333 0.289181
R480 VGND.n489 VGND.n0 0.27022
R481 VGND.n379 VGND.n378 0.2683
R482 VGND.n301 VGND.n141 0.2683
R483 VGND.n186 VGND.n161 0.256021
R484 VGND.n338 VGND.n110 0.250193
R485 VGND.n447 VGND.n444 0.243514
R486 VGND.n333 VGND.n332 0.243383
R487 VGND VGND.n224 0.243171
R488 VGND.n258 VGND.n257 0.241078
R489 VGND.n257 VGND.n256 0.241078
R490 VGND.n17 VGND.n2 0.241078
R491 VGND.n481 VGND.n480 0.241078
R492 VGND.n480 VGND.n479 0.241078
R493 VGND VGND.n224 0.237591
R494 VGND.n405 VGND.n404 0.22226
R495 VGND.n380 VGND.n379 0.221084
R496 VGND.n301 VGND.n300 0.221084
R497 VGND.n332 VGND.n331 0.216589
R498 VGND.n216 VGND.n213 0.208
R499 VGND.n283 VGND.n267 0.201227
R500 VGND.n87 VGND 0.196056
R501 VGND.n381 VGND.n380 0.193014
R502 VGND.n300 VGND.n299 0.193014
R503 VGND.n331 VGND.n330 0.189923
R504 VGND.n247 VGND 0.180825
R505 VGND.n30 VGND 0.180825
R506 VGND.n256 VGND.n255 0.180789
R507 VGND.n487 VGND.n2 0.180789
R508 VGND.n18 VGND.n17 0.180789
R509 VGND.n479 VGND.n478 0.180789
R510 VGND.n237 VGND.n236 0.177986
R511 VGND.n21 VGND.n20 0.177986
R512 VGND.n48 VGND.n47 0.177986
R513 VGND.n330 VGND.n329 0.177878
R514 VGND.n382 VGND.n381 0.172356
R515 VGND.n299 VGND.n298 0.172356
R516 VGND.n186 VGND.n185 0.165165
R517 VGND.n250 VGND.n249 0.163289
R518 VGND.n33 VGND.n32 0.163289
R519 VGND.n329 VGND.n328 0.161737
R520 VGND.n244 VGND.n243 0.159539
R521 VGND.n28 VGND.n27 0.159539
R522 VGND.n57 VGND.n42 0.159539
R523 VGND.n459 VGND.n73 0.158526
R524 VGND.n236 VGND.n220 0.158325
R525 VGND.n20 VGND.n19 0.158325
R526 VGND.n48 VGND.n40 0.158325
R527 VGND.n383 VGND.n382 0.155671
R528 VGND.n298 VGND.n297 0.155671
R529 VGND.n185 VGND.n184 0.152148
R530 VGND.n388 VGND.n387 0.150927
R531 VGND.n328 VGND.n327 0.149148
R532 VGND.n386 VGND.n90 0.149023
R533 VGND.n385 VGND.n91 0.147167
R534 VGND.n295 VGND.n147 0.147167
R535 VGND.n184 VGND.n183 0.145833
R536 VGND.n242 VGND.n240 0.145789
R537 VGND.n26 VGND.n24 0.145789
R538 VGND.n45 VGND.n44 0.145789
R539 VGND.n384 VGND.n92 0.144762
R540 VGND.n296 VGND.n146 0.144762
R541 VGND.n384 VGND.n383 0.143511
R542 VGND.n297 VGND.n296 0.143511
R543 VGND.n150 VGND.n149 0.143335
R544 VGND.n383 VGND.n93 0.14301
R545 VGND.n297 VGND.n145 0.14301
R546 VGND.n327 VGND.n326 0.142866
R547 VGND.n382 VGND.n94 0.1413
R548 VGND.n298 VGND.n144 0.1413
R549 VGND.n381 VGND.n95 0.13963
R550 VGND.n299 VGND.n143 0.13963
R551 VGND.n380 VGND.n96 0.138
R552 VGND.n300 VGND.n142 0.138
R553 VGND.n249 VGND.n247 0.137986
R554 VGND.n32 VGND.n30 0.137986
R555 VGND.n183 VGND.n182 0.136464
R556 VGND.n379 VGND.n97 0.136407
R557 VGND.n302 VGND.n301 0.136407
R558 VGND.n454 VGND.n453 0.134991
R559 VGND.n378 VGND.n98 0.134851
R560 VGND.n303 VGND.n141 0.134851
R561 VGND.n385 VGND.n384 0.134721
R562 VGND.n296 VGND.n295 0.134721
R563 VGND.n326 VGND.n325 0.133592
R564 VGND.n377 VGND.n99 0.13333
R565 VGND.n182 VGND.n181 0.131588
R566 VGND.n239 VGND.n238 0.130789
R567 VGND.n23 VGND.n22 0.130789
R568 VGND.n325 VGND.n324 0.127631
R569 VGND.n348 VGND.n109 0.127631
R570 VGND.n386 VGND.n385 0.127467
R571 VGND.n295 VGND.n294 0.127467
R572 VGND.n181 VGND.n180 0.126098
R573 VGND.n324 VGND.n323 0.123294
R574 VGND.n238 VGND.n237 0.123289
R575 VGND.n22 VGND.n21 0.123289
R576 VGND.n47 VGND.n46 0.123289
R577 VGND.n389 VGND.n388 0.122249
R578 VGND.n352 VGND.n109 0.122221
R579 VGND.n347 VGND.n110 0.122211
R580 VGND.n180 VGND.n179 0.121629
R581 VGND.n387 VGND.n386 0.121573
R582 VGND.n294 VGND.n293 0.121573
R583 VGND.n403 VGND.n46 0.120789
R584 VGND.n174 VGND.n173 0.119457
R585 VGND.n179 VGND.n178 0.118673
R586 VGND.n353 VGND.n352 0.117844
R587 VGND.n174 VGND.n73 0.117211
R588 VGND.n178 VGND.n177 0.114913
R589 VGND.n354 VGND.n353 0.114675
R590 VGND.n177 VGND.n176 0.113743
R591 VGND.n337 VGND.n112 0.112734
R592 VGND.n336 VGND.n335 0.112578
R593 VGND.n253 VGND.n250 0.112039
R594 VGND.n36 VGND.n33 0.112039
R595 VGND.n334 VGND.n113 0.111718
R596 VGND.n333 VGND.n114 0.111507
R597 VGND.n319 VGND.n318 0.111202
R598 VGND.n354 VGND.n107 0.111202
R599 VGND.n294 VGND.n148 0.11115
R600 VGND.n240 VGND.n239 0.110789
R601 VGND.n24 VGND.n23 0.110789
R602 VGND.n402 VGND.n45 0.110789
R603 VGND.n176 VGND.n175 0.110741
R604 VGND.n332 VGND.n115 0.110644
R605 VGND.n175 VGND.n174 0.110231
R606 VGND.n331 VGND.n116 0.110139
R607 VGND.n318 VGND.n317 0.110119
R608 VGND.n330 VGND.n117 0.109632
R609 VGND.n187 VGND.n186 0.109257
R610 VGND.n358 VGND.n107 0.109256
R611 VGND.n329 VGND.n118 0.109053
R612 VGND.n185 VGND.n162 0.10874
R613 VGND.n328 VGND.n119 0.10854
R614 VGND.n184 VGND.n163 0.108513
R615 VGND.n183 VGND.n164 0.108352
R616 VGND.n182 VGND.n165 0.108122
R617 VGND.n327 VGND.n120 0.108023
R618 VGND.n326 VGND.n121 0.107796
R619 VGND.n180 VGND.n167 0.107722
R620 VGND.n181 VGND.n166 0.107592
R621 VGND.n179 VGND.n168 0.107552
R622 VGND.n177 VGND.n170 0.10751
R623 VGND.n325 VGND.n122 0.107273
R624 VGND.n349 VGND.n348 0.107273
R625 VGND.n317 VGND.n316 0.107182
R626 VGND.n304 VGND.n139 0.107096
R627 VGND.n175 VGND.n172 0.107092
R628 VGND.n324 VGND.n123 0.107042
R629 VGND.n350 VGND.n109 0.107042
R630 VGND.n178 VGND.n169 0.10701
R631 VGND.n176 VGND.n171 0.106962
R632 VGND.n323 VGND.n124 0.10687
R633 VGND.n352 VGND.n351 0.10687
R634 VGND.n321 VGND.n126 0.106635
R635 VGND.n353 VGND.n108 0.106635
R636 VGND.n375 VGND.n101 0.106426
R637 VGND.n359 VGND.n358 0.106367
R638 VGND.n319 VGND.n127 0.1061
R639 VGND.n355 VGND.n354 0.1061
R640 VGND.n317 VGND.n129 0.10604
R641 VGND.n358 VGND.n357 0.10604
R642 VGND.n315 VGND.n131 0.105977
R643 VGND.n361 VGND.n360 0.105977
R644 VGND.n310 VGND.n136 0.105973
R645 VGND.n368 VGND.n103 0.105973
R646 VGND.n318 VGND.n128 0.10592
R647 VGND.n356 VGND.n107 0.10592
R648 VGND.n374 VGND.n102 0.105907
R649 VGND.n311 VGND.n135 0.105848
R650 VGND.n367 VGND.n366 0.105848
R651 VGND.n309 VGND.n137 0.10578
R652 VGND.n370 VGND.n369 0.10578
R653 VGND.n314 VGND.n132 0.105731
R654 VGND.n362 VGND.n105 0.105731
R655 VGND.n316 VGND.n315 0.105665
R656 VGND.n312 VGND.n134 0.105663
R657 VGND.n365 VGND.n104 0.105663
R658 VGND.n313 VGND.n133 0.105542
R659 VGND.n364 VGND.n363 0.105542
R660 VGND.n316 VGND.n130 0.105493
R661 VGND.n359 VGND.n106 0.105493
R662 VGND.n360 VGND.n359 0.104886
R663 VGND.n292 VGND.n150 0.104495
R664 VGND.n315 VGND.n314 0.104166
R665 VGND.n360 VGND.n105 0.104166
R666 VGND.n404 uio_out[1] 0.10346
R667 VGND.n313 VGND.n312 0.102551
R668 VGND.n314 VGND.n313 0.102053
R669 VGND.n364 VGND.n105 0.102053
R670 VGND.n320 VGND.n319 0.101891
R671 VGND.n365 VGND.n364 0.101858
R672 VGND.n312 VGND.n311 0.101493
R673 VGND.n366 VGND.n365 0.101493
R674 VGND.n311 VGND.n310 0.100967
R675 VGND.n366 VGND.n103 0.100967
R676 VGND.n308 VGND.n307 0.100958
R677 VGND.n309 VGND.n308 0.100445
R678 VGND.n375 VGND.n374 0.100376
R679 VGND.n310 VGND.n309 0.100187
R680 VGND.n370 VGND.n103 0.100187
R681 VGND.n73 VGND.n72 0.0973571
R682 VGND.n244 VGND.n242 0.095789
R683 VGND.n28 VGND.n26 0.095789
R684 VGND.n44 VGND.n42 0.095789
R685 VGND.n453 VGND.n452 0.0954338
R686 VGND.n448 VGND.n85 0.0928432
R687 VGND.n323 VGND.n322 0.0895217
R688 VGND.n457 VGND.n456 0.0873393
R689 VGND.n387 VGND.n89 0.085643
R690 VGND.n204 VGND 0.0854123
R691 VGND.n255 VGND.n220 0.083
R692 VGND.n19 VGND.n18 0.083
R693 VGND.n478 VGND.n40 0.083
R694 VGND.n308 VGND.n138 0.0814084
R695 VGND.n376 VGND.n100 0.0802603
R696 VGND.n101 VGND.n100 0.0782828
R697 VGND.n488 VGND.n487 0.078
R698 VGND.n388 VGND.n90 0.0779701
R699 VGND.n374 VGND.n373 0.0771258
R700 VGND.n348 VGND.n347 0.0762778
R701 VGND.n452 VGND.n451 0.0754235
R702 VGND.n91 VGND.n90 0.0751329
R703 VGND.n448 VGND.n447 0.0739655
R704 VGND.n148 VGND.n147 0.0735315
R705 VGND.n92 VGND.n91 0.0731
R706 VGND.n147 VGND.n146 0.0731
R707 VGND.n456 VGND.n79 0.0724725
R708 VGND.n93 VGND.n92 0.0701066
R709 VGND.n146 VGND.n145 0.0701066
R710 VGND.n94 VGND.n93 0.067836
R711 VGND.n145 VGND.n144 0.067836
R712 VGND.n307 VGND.n306 0.0669444
R713 VGND.n95 VGND.n94 0.06562
R714 VGND.n144 VGND.n143 0.06562
R715 VGND.t55 VGND.n210 0.0650946
R716 VGND.t7 VGND.n246 0.0650946
R717 VGND.t7 VGND.n222 0.0650946
R718 VGND.t79 VGND.n10 0.0650946
R719 VGND.n96 VGND.n95 0.0634565
R720 VGND.n143 VGND.n142 0.0634565
R721 VGND.n451 VGND.n450 0.0614573
R722 VGND.n285 VGND 0.061
R723 VGND.n265 VGND 0.061
R724 VGND.n391 VGND 0.061
R725 VGND.n77 VGND 0.061
R726 VGND.n76 VGND 0.061
R727 VGND.n461 VGND 0.061
R728 VGND.n189 VGND 0.061
R729 VGND.n159 VGND 0.061
R730 VGND.n446 VGND 0.061
R731 VGND.n88 VGND 0.061
R732 VGND.n97 VGND.n96 0.061
R733 VGND.n140 VGND 0.061
R734 VGND.n291 VGND 0.061
R735 VGND.n275 VGND 0.061
R736 VGND.n269 VGND 0.061
R737 VGND.n302 VGND.n142 0.061
R738 VGND.n340 VGND 0.061
R739 VGND.n346 VGND 0.061
R740 VGND.n372 VGND 0.061
R741 VGND.n193 VGND 0.061
R742 VGND.n282 VGND 0.061
R743 VGND.n81 VGND.n80 0.0607651
R744 VGND.n227 VGND 0.0605
R745 VGND VGND.n13 0.0605
R746 VGND.n58 VGND 0.0605
R747 VGND.n389 VGND.n89 0.060354
R748 VGND.n98 VGND.n97 0.0589402
R749 VGND.n303 VGND.n302 0.0589402
R750 VGND.n450 VGND.n449 0.0585315
R751 VGND.n293 VGND.n149 0.0568276
R752 VGND.n99 VGND.n98 0.0565916
R753 VGND.n304 VGND.n303 0.0565916
R754 uo_out[4] VGND.n489 0.0555
R755 VGND.n85 VGND.n84 0.0547113
R756 VGND.n100 VGND.n99 0.0546283
R757 VGND.n454 VGND.n81 0.0545351
R758 VGND.n456 VGND.n455 0.0537058
R759 VGND.n138 VGND.n137 0.0535756
R760 VGND.n376 VGND.n375 0.0505564
R761 VGND.n102 VGND.n101 0.0497148
R762 VGND.n84 VGND.n83 0.0483673
R763 VGND.n305 VGND.n304 0.048347
R764 VGND.n369 VGND.n102 0.0478846
R765 VGND.n137 VGND.n136 0.04594
R766 VGND.n369 VGND.n368 0.04594
R767 VGND VGND.n87 0.0445
R768 VGND.n136 VGND.n135 0.0440235
R769 VGND.n368 VGND.n367 0.0440235
R770 VGND.n488 VGND.n1 0.043
R771 VGND.n135 VGND.n134 0.0421344
R772 VGND.n367 VGND.n104 0.0421344
R773 VGND.n83 VGND.n82 0.0419304
R774 VGND.n173 VGND.n72 0.0411957
R775 VGND.n307 VGND.n139 0.0409767
R776 VGND.n134 VGND.n133 0.0401312
R777 VGND.n363 VGND.n104 0.0401312
R778 VGND.n149 VGND.n148 0.0397586
R779 VGND.n133 VGND.n132 0.0386127
R780 VGND.n363 VGND.n362 0.0386127
R781 VGND.n306 VGND.n305 0.0384989
R782 VGND.n132 VGND.n131 0.0365
R783 VGND.n362 VGND.n361 0.0365
R784 VGND.n460 VGND.n72 0.0356429
R785 VGND.n173 VGND.n172 0.0355141
R786 VGND.n131 VGND.n130 0.0351481
R787 VGND.n361 VGND.n106 0.0351481
R788 VGND.n172 VGND.n171 0.0337308
R789 VGND.n130 VGND.n129 0.0332724
R790 VGND.n357 VGND.n106 0.0332724
R791 VGND.n338 VGND.n337 0.032543
R792 VGND.n444 VGND.n393 0.0319281
R793 VGND.n171 VGND.n170 0.0317753
R794 VGND.n129 VGND.n128 0.0313454
R795 VGND.n357 VGND.n356 0.0313454
R796 VGND.n349 VGND.n110 0.0307408
R797 VGND.n170 VGND.n169 0.0302379
R798 VGND.n128 VGND.n127 0.0299334
R799 VGND.n356 VGND.n355 0.0299334
R800 VGND.n322 VGND.n321 0.0298333
R801 VGND.n169 VGND.n168 0.0283213
R802 VGND.n127 VGND.n126 0.0279441
R803 VGND.n355 VGND.n108 0.0279441
R804 VGND.n80 VGND.n79 0.0273067
R805 VGND.n168 VGND.n167 0.0266297
R806 VGND.n126 VGND.n124 0.0263649
R807 VGND.n351 VGND.n108 0.0263649
R808 VGND.n139 VGND.n138 0.0255726
R809 VGND.n167 VGND.n166 0.024961
R810 VGND.n441 VGND.n394 0.0249162
R811 VGND.n430 VGND.n423 0.0249162
R812 VGND.n124 VGND.n123 0.0247963
R813 VGND.n351 VGND.n350 0.0247963
R814 VGND.n166 VGND.n165 0.0233919
R815 VGND.n373 VGND.n370 0.02322
R816 VGND.n123 VGND.n122 0.0231622
R817 VGND.n350 VGND.n349 0.0231622
R818 VGND.n165 VGND.n164 0.0218333
R819 VGND.n243 VGND.n227 0.02175
R820 VGND.n27 VGND.n13 0.02175
R821 VGND.n58 VGND.n57 0.02175
R822 VGND.n443 VGND.n442 0.02162
R823 VGND.n424 VGND.n86 0.02162
R824 VGND.n122 VGND.n121 0.02162
R825 VGND.n460 VGND.n459 0.0212439
R826 VGND.n293 VGND.n292 0.0200345
R827 VGND.n164 VGND.n163 0.0199247
R828 VGND.n121 VGND.n120 0.0197957
R829 VGND.n163 VGND.n162 0.0186867
R830 VGND.n120 VGND.n119 0.0185662
R831 VGND.n455 VGND.n454 0.0170759
R832 VGND.n187 VGND.n162 0.0168721
R833 VGND.n119 VGND.n118 0.016764
R834 VGND.n0 uo_out[5] 0.0157601
R835 VGND.n398 uo_out[6] 0.0157601
R836 VGND.n399 uo_out[7] 0.0157601
R837 VGND.n400 uio_out[0] 0.0157601
R838 VGND.n401 uio_out[1] 0.0157601
R839 VGND.n405 uio_out[2] 0.0157601
R840 VGND.n406 uio_out[3] 0.0157601
R841 VGND.n407 uio_out[4] 0.0157601
R842 VGND.n408 uio_out[5] 0.0157601
R843 VGND.n409 uio_out[6] 0.0157601
R844 VGND.n410 uio_out[7] 0.0157601
R845 VGND.n411 uio_oe[0] 0.0157601
R846 VGND.n412 uio_oe[1] 0.0157601
R847 VGND.n413 uio_oe[2] 0.0157601
R848 VGND.n414 uio_oe[3] 0.0157601
R849 VGND.n415 uio_oe[4] 0.0157601
R850 VGND.n416 uio_oe[5] 0.0157601
R851 VGND.n417 uio_oe[6] 0.0157601
R852 VGND.n418 uio_oe[7] 0.0157601
R853 VGND.n79 VGND.n78 0.0153179
R854 VGND.n188 VGND.n187 0.0150695
R855 VGND.n118 VGND.n117 0.0149737
R856 VGND.n117 VGND.n116 0.0138158
R857 uo_out[5] VGND.n0 0.0137
R858 uo_out[6] VGND.n398 0.0137
R859 uo_out[7] VGND.n399 0.0137
R860 uio_out[0] VGND.n400 0.0137
R861 uio_out[1] VGND.n401 0.0137
R862 uio_out[2] VGND.n405 0.0137
R863 uio_out[3] VGND.n406 0.0137
R864 uio_out[4] VGND.n407 0.0137
R865 uio_out[5] VGND.n408 0.0137
R866 uio_out[6] VGND.n409 0.0137
R867 uio_out[7] VGND.n410 0.0137
R868 uio_oe[0] VGND.n411 0.0137
R869 uio_oe[1] VGND.n412 0.0137
R870 uio_oe[2] VGND.n413 0.0137
R871 uio_oe[3] VGND.n414 0.0137
R872 uio_oe[4] VGND.n415 0.0137
R873 uio_oe[5] VGND.n416 0.0137
R874 uio_oe[6] VGND.n417 0.0137
R875 uio_oe[7] VGND.n418 0.0137
R876 VGND.n321 VGND.n320 0.0132838
R877 VGND.n439 VGND.n395 0.0131992
R878 VGND.n433 VGND.n425 0.0131992
R879 VGND.n441 VGND.n396 0.0131916
R880 VGND.n426 VGND.n423 0.0131916
R881 VGND.n426 VGND.n421 0.0131916
R882 VGND.n419 VGND.n396 0.0131916
R883 VGND.n419 VGND.n395 0.0130858
R884 VGND.n425 VGND.n421 0.0130858
R885 VGND.n82 VGND.n81 0.0121797
R886 VGND.n116 VGND.n115 0.012041
R887 VGND.n440 VGND.n420 0.0115476
R888 VGND.n437 VGND.n435 0.0115476
R889 VGND.n434 VGND.n422 0.0115476
R890 VGND.n431 VGND.n427 0.0115476
R891 VGND.n428 VGND.n422 0.0115476
R892 VGND.n432 VGND.n431 0.0115476
R893 VGND.n436 VGND.n420 0.0115476
R894 VGND.n438 VGND.n437 0.0115476
R895 VGND.n438 VGND.n397 0.0115476
R896 VGND.n432 VGND.n429 0.0115476
R897 VGND.n429 VGND.n428 0.0115476
R898 VGND.n436 VGND.n397 0.0115476
R899 VGND.n115 VGND.n114 0.0105654
R900 VGND.n403 VGND.n402 0.0105
R901 VGND.n457 VGND.n78 0.00934499
R902 VGND.n449 VGND.n448 0.00920833
R903 VGND.n114 VGND.n113 0.00883987
R904 VGND.n453 VGND.n82 0.00874622
R905 VGND.n452 VGND.n83 0.0077971
R906 VGND.n336 VGND.n113 0.00737948
R907 VGND.n451 VGND.n84 0.00643951
R908 VGND.n337 VGND.n336 0.00594625
R909 VGND.n188 VGND.n161 0.00588981
R910 VGND.n455 VGND.n80 0.00446192
R911 VGND.n450 VGND.n85 0.00434654
R912 VGND.n235 VGND.n219 0.00166667
R913 VGND.n483 VGND.n7 0.00166667
R914 VGND.n49 VGND.n39 0.00166667
R915 VGND.t7 VGND.n235 0.00133332
R916 VGND.n483 VGND.t79 0.00133332
R917 VGND.n477 VGND.n49 0.00133332
R918 VGND.n217 VGND.n208 0.001
R919 VGND.n232 VGND.n217 0.001
R920 VGND.n233 VGND.n218 0.001
R921 VGND.n486 VGND.n3 0.001
R922 VGND.n486 VGND.n485 0.001
R923 VGND.n6 VGND.n4 0.001
R924 VGND.n37 VGND.n8 0.001
R925 VGND.n50 VGND.n37 0.001
R926 VGND.n51 VGND.n38 0.001
R927 VGND.t55 VGND.n208 0.001
R928 VGND.n232 VGND.n218 0.001
R929 VGND.n233 VGND.n219 0.001
R930 VGND.t7 VGND.n3 0.001
R931 VGND.n485 VGND.n4 0.001
R932 VGND.n7 VGND.n6 0.001
R933 VGND.t79 VGND.n8 0.001
R934 VGND.n50 VGND.n38 0.001
R935 VGND.n51 VGND.n39 0.001
R936 uo_out[1].n3 uo_out[1].t2 15.0005
R937 uo_out[1] uo_out[1].n3 13.4668
R938 uo_out[1].n2 uo_out[1].n1 9.01747
R939 uo_out[1].n2 uo_out[1] 8.9065
R940 uo_out[1].n0 uo_out[1].t1 8.53421
R941 uo_out[1].n0 uo_out[1].t0 6.13626
R942 uo_out[1].n1 uo_out[1].n0 0.100612
R943 uo_out[1].n1 uo_out[1] 0.0585899
R944 uo_out[1].n3 uo_out[1] 0.04098
R945 uo_out[1] uo_out[1].n2 0.00678571
R946 VDPWR.n7 VDPWR.t1 34.1026
R947 VDPWR.n5 VDPWR.t17 34.1026
R948 VDPWR.n80 VDPWR.t46 34.1026
R949 VDPWR.n79 VDPWR.t3 34.1026
R950 VDPWR.n77 VDPWR.t52 34.1026
R951 VDPWR.n76 VDPWR.t40 34.1026
R952 VDPWR.n35 VDPWR.t62 34.1026
R953 VDPWR.n33 VDPWR.t49 34.1026
R954 VDPWR.n31 VDPWR.t32 34.1026
R955 VDPWR.n24 VDPWR.t24 34.1026
R956 VDPWR.n150 VDPWR.t8 34.1026
R957 VDPWR.n163 VDPWR.t57 34.1026
R958 VDPWR.n161 VDPWR.t66 34.1026
R959 VDPWR.n54 VDPWR.t83 34.1026
R960 VDPWR.n75 VDPWR.t87 34.1026
R961 VDPWR.n78 VDPWR.t38 34.1026
R962 VDPWR.n81 VDPWR.t26 34.1026
R963 VDPWR.n82 VDPWR.t28 34.1026
R964 VDPWR.n83 VDPWR.t59 34.1026
R965 VDPWR.n84 VDPWR.t72 34.1026
R966 VDPWR.n0 VDPWR.t6 34.1026
R967 VDPWR.n230 VDPWR.n173 19.7403
R968 VDPWR VDPWR.n7 18.2059
R969 VDPWR VDPWR.n5 18.2059
R970 VDPWR VDPWR.n80 18.2059
R971 VDPWR VDPWR.n79 18.2059
R972 VDPWR VDPWR.n77 18.2059
R973 VDPWR VDPWR.n76 18.2059
R974 VDPWR VDPWR.n35 18.2059
R975 VDPWR VDPWR.n33 18.2059
R976 VDPWR VDPWR.n31 18.2059
R977 VDPWR VDPWR.n24 18.2059
R978 VDPWR VDPWR.n150 18.2059
R979 VDPWR VDPWR.n163 18.2059
R980 VDPWR VDPWR.n161 18.2059
R981 VDPWR VDPWR.n54 18.2059
R982 VDPWR VDPWR.n75 18.2059
R983 VDPWR VDPWR.n78 18.2059
R984 VDPWR VDPWR.n81 18.2059
R985 VDPWR VDPWR.n82 18.2059
R986 VDPWR VDPWR.n83 18.2059
R987 VDPWR VDPWR.n84 18.2059
R988 VDPWR VDPWR.n0 18.2059
R989 VDPWR.n230 VDPWR.n229 18.0005
R990 VDPWR.n220 VDPWR.t51 17.378
R991 VDPWR.n207 VDPWR.t20 17.378
R992 VDPWR.n190 VDPWR.t35 17.378
R993 VDPWR.n221 VDPWR.t48 17.3693
R994 VDPWR.n205 VDPWR.t36 17.3693
R995 VDPWR.n189 VDPWR.t5 17.3693
R996 VDPWR.n7 VDPWR.t2 17.0233
R997 VDPWR.n5 VDPWR.t18 17.0233
R998 VDPWR.n80 VDPWR.t47 17.0233
R999 VDPWR.n79 VDPWR.t4 17.0233
R1000 VDPWR.n77 VDPWR.t53 17.0233
R1001 VDPWR.n76 VDPWR.t41 17.0233
R1002 VDPWR.n35 VDPWR.t63 17.0233
R1003 VDPWR.n33 VDPWR.t50 17.0233
R1004 VDPWR.n31 VDPWR.t33 17.0233
R1005 VDPWR.n24 VDPWR.t25 17.0233
R1006 VDPWR.n150 VDPWR.t9 17.0233
R1007 VDPWR.n163 VDPWR.t58 17.0233
R1008 VDPWR.n161 VDPWR.t67 17.0233
R1009 VDPWR.n54 VDPWR.t84 17.0233
R1010 VDPWR.n75 VDPWR.t88 17.0233
R1011 VDPWR.n78 VDPWR.t39 17.0233
R1012 VDPWR.n81 VDPWR.t27 17.0233
R1013 VDPWR.n82 VDPWR.t29 17.0233
R1014 VDPWR.n83 VDPWR.t60 17.0233
R1015 VDPWR.n84 VDPWR.t73 17.0233
R1016 VDPWR.n0 VDPWR.t7 17.0233
R1017 VDPWR.n220 VDPWR.t15 17.0005
R1018 VDPWR.t10 VDPWR.n188 17.0005
R1019 VDPWR.n227 VDPWR.t10 17.0005
R1020 VDPWR.n207 VDPWR.t16 17.0005
R1021 VDPWR.t23 VDPWR.n209 17.0005
R1022 VDPWR.t23 VDPWR.n211 17.0005
R1023 VDPWR.t23 VDPWR.n200 17.0005
R1024 VDPWR.n190 VDPWR.t19 17.0005
R1025 VDPWR.t10 VDPWR.n174 17.0005
R1026 VDPWR.t10 VDPWR.n181 17.0005
R1027 VDPWR.t10 VDPWR.n194 17.0005
R1028 VDPWR.n223 VDPWR.t23 17.0005
R1029 VDPWR.n231 VDPWR.n230 12.4694
R1030 VDPWR.n171 VDPWR.n170 9.2117
R1031 VDPWR.n167 VDPWR.n153 9.18823
R1032 VDPWR.n171 VDPWR.n18 9.18823
R1033 VDPWR.n171 VDPWR.n17 9.05079
R1034 VDPWR.n168 VDPWR.n167 9.0005
R1035 VDPWR.n169 VDPWR.n18 9.0005
R1036 VDPWR.n168 VDPWR.n21 9.0005
R1037 VDPWR.n169 VDPWR.n17 9.0005
R1038 VDPWR.n168 VDPWR.n19 9.0005
R1039 VDPWR.n170 VDPWR.n169 9.0005
R1040 VDPWR.n157 VDPWR.n156 9.0005
R1041 VDPWR.n154 VDPWR.n11 9.0005
R1042 VDPWR.n235 VDPWR.n13 9.0005
R1043 VDPWR.n218 VDPWR.t13 8.80285
R1044 VDPWR.n196 VDPWR.t69 8.80285
R1045 VDPWR.n184 VDPWR.t44 8.80285
R1046 VDPWR.t0 VDPWR.n201 8.501
R1047 VDPWR.t23 VDPWR.n215 8.47111
R1048 VDPWR.t23 VDPWR.n217 8.47111
R1049 VDPWR.t10 VDPWR.n185 8.47111
R1050 VDPWR.t10 VDPWR.n178 8.47111
R1051 VDPWR.t10 VDPWR.n176 8.47111
R1052 VDPWR.n225 VDPWR.n197 8.47111
R1053 VDPWR.n224 VDPWR.n198 8.47111
R1054 VDPWR.n183 VDPWR.t42 6.07323
R1055 VDPWR.n216 VDPWR.t11 6.073
R1056 VDPWR.n177 VDPWR.t68 6.073
R1057 VDPWR.n88 VDPWR.n87 6.01045
R1058 VDPWR.n187 VDPWR.t55 5.98925
R1059 VDPWR.n175 VDPWR.t54 5.98882
R1060 VDPWR.n214 VDPWR.t22 5.98825
R1061 VDPWR.n212 VDPWR.t21 5.98825
R1062 VDPWR.n179 VDPWR.t30 5.98825
R1063 VDPWR.n193 VDPWR.t31 5.98825
R1064 VDPWR.n6 VDPWR 5.96901
R1065 VDPWR.n151 VDPWR.n149 5.84778
R1066 VDPWR.t10 VDPWR.n186 5.61485
R1067 VDPWR.t23 VDPWR.n213 5.61485
R1068 VDPWR.t10 VDPWR.n180 5.61485
R1069 VDPWR.t10 VDPWR.n226 5.61485
R1070 VDPWR.n232 VDPWR 5.2541
R1071 VDPWR.n93 VDPWR.n92 5.21746
R1072 VDPWR VDPWR.n250 4.73
R1073 VDPWR.n239 VDPWR 4.6152
R1074 VDPWR.n153 VDPWR.n152 4.53071
R1075 VDPWR.n166 VDPWR.n22 4.51901
R1076 VDPWR.n165 VDPWR.n16 4.50989
R1077 VDPWR.n85 VDPWR 4.13588
R1078 VDPWR.n86 VDPWR 3.92388
R1079 VDPWR.n88 VDPWR 3.88095
R1080 VDPWR.n87 VDPWR 3.84419
R1081 VDPWR.n162 VDPWR 3.66357
R1082 VDPWR.n89 VDPWR 3.41222
R1083 VDPWR.t23 VDPWR.n210 3.33162
R1084 VDPWR.t10 VDPWR.n192 3.30723
R1085 VDPWR.t23 VDPWR.n206 3.30706
R1086 VDPWR.n164 VDPWR 3.28289
R1087 VDPWR.n156 VDPWR.n155 3.0005
R1088 VDPWR.n11 VDPWR.n9 3.0005
R1089 VDPWR.n236 VDPWR.n235 3.0005
R1090 VDPWR.n151 VDPWR 2.98934
R1091 VDPWR.t23 VDPWR.n222 2.72512
R1092 VDPWR.n239 VDPWR.n238 2.5318
R1093 VDPWR.n25 VDPWR 2.53128
R1094 VDPWR.n136 VDPWR.n34 2.46388
R1095 VDPWR.t23 VDPWR.n204 2.29759
R1096 VDPWR.n153 VDPWR.n20 2.27162
R1097 VDPWR.n159 VDPWR.n12 2.26628
R1098 VDPWR.n172 VDPWR.n171 2.2505
R1099 VDPWR.n168 VDPWR.n20 2.2505
R1100 VDPWR.n169 VDPWR.n15 2.2505
R1101 VDPWR.n233 VDPWR.n12 2.2505
R1102 VDPWR.n235 VDPWR.n234 2.2505
R1103 VDPWR.n90 VDPWR 2.15229
R1104 VDPWR.n203 VDPWR 2.0605
R1105 VDPWR.n32 VDPWR 1.94477
R1106 VDPWR.n232 VDPWR.n231 1.89976
R1107 VDPWR.n91 VDPWR 1.74056
R1108 VDPWR.n93 VDPWR 1.53994
R1109 VDPWR.n199 VDPWR 1.53643
R1110 VDPWR.n233 VDPWR.n232 1.47736
R1111 VDPWR.n231 VDPWR.n172 1.46416
R1112 VDPWR.n92 VDPWR 1.39911
R1113 VDPWR.n95 VDPWR 1.19117
R1114 VDPWR.n137 VDPWR 1.1824
R1115 VDPWR.n234 VDPWR.n14 1.14638
R1116 VDPWR.n90 VDPWR.n89 1.035
R1117 VDPWR.n94 VDPWR.n93 0.923201
R1118 VDPWR.n116 VDPWR 0.895684
R1119 VDPWR.n135 VDPWR 0.886
R1120 VDPWR.n184 VDPWR.n182 0.854038
R1121 VDPWR.n219 VDPWR.n218 0.851125
R1122 VDPWR.n221 VDPWR.n219 0.805789
R1123 VDPWR.n189 VDPWR.n182 0.803932
R1124 VDPWR.t10 VDPWR.n182 0.802654
R1125 VDPWR.t23 VDPWR.n219 0.800901
R1126 VDPWR.n138 VDPWR.n137 0.767737
R1127 VDPWR.n85 VDPWR.n1 0.762233
R1128 VDPWR.n228 VDPWR 0.543
R1129 VDPWR.n144 VDPWR.n23 0.531002
R1130 VDPWR.n61 VDPWR.n60 0.507992
R1131 VDPWR.n222 VDPWR.n220 0.410237
R1132 VDPWR.t0 VDPWR.n195 0.40574
R1133 VDPWR.n91 VDPWR.n90 0.393052
R1134 VDPWR.n204 VDPWR.n203 0.392162
R1135 VDPWR.n222 VDPWR.n221 0.389189
R1136 VDPWR.n205 VDPWR.n204 0.374189
R1137 VDPWR.n87 VDPWR.n86 0.363276
R1138 VDPWR.n202 VDPWR.t0 0.341
R1139 VDPWR.n192 VDPWR.n189 0.336433
R1140 VDPWR.n206 VDPWR.n205 0.336118
R1141 VDPWR.n164 VDPWR.n162 0.334929
R1142 VDPWR.n92 VDPWR.n91 0.332665
R1143 VDPWR.n208 VDPWR.n206 0.331746
R1144 VDPWR.n192 VDPWR.n191 0.331445
R1145 VDPWR.n36 VDPWR.n34 0.330588
R1146 VDPWR.n89 VDPWR.n88 0.323555
R1147 VDPWR.n165 VDPWR.n164 0.312824
R1148 VDPWR.n137 VDPWR.n136 0.305164
R1149 VDPWR.n226 VDPWR.n225 0.300775
R1150 VDPWR.n86 VDPWR.n85 0.289257
R1151 VDPWR.n62 VDPWR.n61 0.2887
R1152 VDPWR.n37 VDPWR.n36 0.280623
R1153 VDPWR.n210 VDPWR 0.273551
R1154 VDPWR.n143 VDPWR.n26 0.251853
R1155 VDPWR.n142 VDPWR.n27 0.2469
R1156 VDPWR.n141 VDPWR.n28 0.24161
R1157 VDPWR.n96 VDPWR.n74 0.24161
R1158 VDPWR.n225 VDPWR.n224 0.241078
R1159 VDPWR.n38 VDPWR.n37 0.240286
R1160 VDPWR.n140 VDPWR.n29 0.237849
R1161 VDPWR.n97 VDPWR.n73 0.237849
R1162 VDPWR.n139 VDPWR.n30 0.234669
R1163 VDPWR.n98 VDPWR.n72 0.234669
R1164 VDPWR.n99 VDPWR.n71 0.231561
R1165 VDPWR.n148 VDPWR.n147 0.230306
R1166 VDPWR.n100 VDPWR.n70 0.226786
R1167 VDPWR.n63 VDPWR.n62 0.225081
R1168 VDPWR.n101 VDPWR.n69 0.22337
R1169 VDPWR.n102 VDPWR.n68 0.219324
R1170 VDPWR.n103 VDPWR.n67 0.217223
R1171 VDPWR.n104 VDPWR.n66 0.213359
R1172 VDPWR.n145 VDPWR.n144 0.212767
R1173 VDPWR.n170 VDPWR.n19 0.2117
R1174 VDPWR.n105 VDPWR.n65 0.211333
R1175 VDPWR.n106 VDPWR.n64 0.208253
R1176 VDPWR VDPWR.n210 0.205841
R1177 VDPWR.n39 VDPWR.n38 0.204702
R1178 VDPWR.n107 VDPWR.n63 0.204642
R1179 VDPWR.n108 VDPWR.n62 0.202722
R1180 VDPWR.n149 VDPWR.n23 0.201278
R1181 VDPWR.n109 VDPWR.n61 0.19982
R1182 VDPWR.n40 VDPWR.n39 0.187779
R1183 VDPWR.n226 VDPWR.n196 0.185825
R1184 VDPWR.n224 VDPWR.n223 0.180789
R1185 VDPWR.n64 VDPWR.n63 0.177266
R1186 VDPWR.n139 VDPWR.n138 0.175862
R1187 VDPWR.n41 VDPWR.n40 0.175509
R1188 VDPWR.n111 VDPWR.n59 0.173049
R1189 VDPWR.n112 VDPWR.n58 0.172207
R1190 VDPWR.n215 VDPWR.n214 0.172039
R1191 VDPWR.n179 VDPWR.n178 0.172039
R1192 VDPWR.n113 VDPWR.n57 0.171374
R1193 VDPWR.n114 VDPWR.n56 0.169731
R1194 VDPWR.n115 VDPWR.n55 0.168921
R1195 VDPWR.n248 VDPWR.n1 0.167396
R1196 VDPWR.n116 VDPWR.n53 0.167325
R1197 VDPWR.n117 VDPWR.n52 0.166538
R1198 VDPWR.n118 VDPWR.n51 0.165758
R1199 VDPWR.n94 VDPWR.n74 0.165337
R1200 VDPWR.n119 VDPWR.n50 0.164986
R1201 VDPWR.n120 VDPWR.n49 0.164221
R1202 VDPWR.n121 VDPWR.n48 0.163463
R1203 VDPWR.n147 VDPWR.n146 0.162204
R1204 VDPWR.n123 VDPWR.n46 0.161968
R1205 VDPWR.n122 VDPWR.n47 0.161968
R1206 VDPWR.n125 VDPWR.n44 0.161231
R1207 VDPWR.n124 VDPWR.n45 0.161231
R1208 VDPWR.n128 VDPWR.n41 0.159776
R1209 VDPWR.n127 VDPWR.n42 0.159776
R1210 VDPWR.n126 VDPWR.n43 0.159776
R1211 VDPWR.n130 VDPWR.n39 0.159059
R1212 VDPWR.n129 VDPWR.n40 0.159059
R1213 VDPWR.n133 VDPWR.n36 0.158348
R1214 VDPWR.n132 VDPWR.n37 0.158348
R1215 VDPWR.n131 VDPWR.n38 0.158348
R1216 VDPWR.n160 VDPWR.n158 0.158044
R1217 VDPWR.n42 VDPWR.n41 0.157911
R1218 VDPWR.n65 VDPWR.n64 0.157621
R1219 VDPWR.n134 VDPWR.n34 0.154546
R1220 VDPWR.n110 VDPWR.n60 0.15242
R1221 VDPWR.n241 VDPWR.n240 0.152188
R1222 VDPWR.n43 VDPWR.n42 0.147308
R1223 VDPWR.n166 VDPWR.n18 0.147167
R1224 VDPWR.n44 VDPWR.n43 0.14126
R1225 VDPWR.n66 VDPWR.n65 0.141098
R1226 VDPWR.n217 VDPWR.n216 0.140789
R1227 VDPWR.n177 VDPWR.n176 0.140789
R1228 VDPWR.n185 VDPWR.n183 0.140789
R1229 VDPWR.n208 VDPWR.n207 0.136382
R1230 VDPWR.n191 VDPWR.n190 0.136382
R1231 VDPWR.n247 VDPWR.n2 0.135022
R1232 VDPWR.n45 VDPWR.n44 0.133682
R1233 VDPWR.n186 VDPWR.n175 0.129236
R1234 VDPWR.n214 VDPWR.n213 0.129236
R1235 VDPWR.n180 VDPWR.n179 0.129236
R1236 VDPWR.n187 VDPWR.n186 0.128325
R1237 VDPWR.n213 VDPWR.n212 0.128325
R1238 VDPWR.n193 VDPWR.n180 0.128325
R1239 VDPWR.n46 VDPWR.n45 0.127233
R1240 VDPWR.n145 VDPWR.n26 0.1269
R1241 VDPWR.n67 VDPWR.n66 0.126475
R1242 VDPWR.n47 VDPWR.n46 0.123269
R1243 VDPWR.n48 VDPWR.n47 0.121562
R1244 VDPWR.n152 VDPWR.n19 0.1171
R1245 VDPWR.n49 VDPWR.n48 0.116891
R1246 VDPWR.n68 VDPWR.n67 0.116337
R1247 VDPWR.n218 VDPWR.n217 0.115789
R1248 VDPWR.n196 VDPWR.n176 0.115789
R1249 VDPWR.n185 VDPWR.n184 0.115789
R1250 VDPWR.n50 VDPWR.n49 0.114401
R1251 VDPWR.n188 VDPWR.n187 0.113
R1252 VDPWR.n212 VDPWR.n211 0.113
R1253 VDPWR.n194 VDPWR.n193 0.113
R1254 VDPWR.n227 VDPWR.n175 0.11175
R1255 VDPWR.n51 VDPWR.n50 0.111106
R1256 VDPWR.n52 VDPWR.n51 0.110556
R1257 VDPWR.n53 VDPWR.n52 0.108981
R1258 VDPWR.n55 VDPWR.n53 0.108669
R1259 VDPWR.n56 VDPWR.n55 0.108583
R1260 VDPWR.n69 VDPWR.n68 0.108277
R1261 VDPWR.n57 VDPWR.n56 0.108072
R1262 VDPWR.n59 VDPWR.n58 0.107345
R1263 VDPWR.n58 VDPWR.n57 0.107234
R1264 VDPWR.n70 VDPWR.n69 0.103826
R1265 VDPWR.n216 VDPWR.n215 0.100789
R1266 VDPWR.n178 VDPWR.n177 0.100789
R1267 VDPWR.n71 VDPWR.n70 0.0994295
R1268 VDPWR.n72 VDPWR.n71 0.096586
R1269 VDPWR.n243 VDPWR.n4 0.0942964
R1270 VDPWR.n140 VDPWR.n139 0.0929227
R1271 VDPWR.n73 VDPWR.n72 0.0929227
R1272 VDPWR.n250 VDPWR.n1 0.0929187
R1273 VDPWR.n141 VDPWR.n140 0.0912154
R1274 VDPWR.n74 VDPWR.n73 0.0912154
R1275 VDPWR.n247 VDPWR.n246 0.0893224
R1276 VDPWR.n142 VDPWR.n141 0.0884738
R1277 VDPWR.n229 VDPWR.n228 0.088
R1278 VDPWR.n143 VDPWR.n142 0.0871337
R1279 VDPWR.n144 VDPWR.n143 0.0864426
R1280 VDPWR.n250 VDPWR.n249 0.0849682
R1281 VDPWR.n27 VDPWR.n26 0.0816497
R1282 VDPWR.n146 VDPWR.n145 0.0787288
R1283 VDPWR.n28 VDPWR.n27 0.0781471
R1284 VDPWR.n96 VDPWR.n95 0.0781471
R1285 VDPWR.n249 VDPWR.n2 0.0761377
R1286 VDPWR.n29 VDPWR.n28 0.0757832
R1287 VDPWR.n97 VDPWR.n96 0.0757832
R1288 VDPWR.n30 VDPWR.n29 0.0734143
R1289 VDPWR.n98 VDPWR.n97 0.0734143
R1290 VDPWR.n245 VDPWR.n2 0.0722058
R1291 VDPWR.n199 VDPWR.n173 0.0717963
R1292 VDPWR.n242 VDPWR.n6 0.071653
R1293 VDPWR.n32 VDPWR.n30 0.071596
R1294 VDPWR.n99 VDPWR.n98 0.071596
R1295 VDPWR.n100 VDPWR.n99 0.0688352
R1296 VDPWR.n111 VDPWR.n110 0.0683607
R1297 VDPWR.n243 VDPWR.n242 0.0679195
R1298 VDPWR.n101 VDPWR.n100 0.0662582
R1299 VDPWR.n203 VDPWR.n200 0.0656852
R1300 VDPWR.n147 VDPWR.n23 0.0656852
R1301 VDPWR.n102 VDPWR.n101 0.0641087
R1302 VDPWR.n95 VDPWR.n94 0.0637952
R1303 VDPWR.n155 VDPWR.n8 0.0627642
R1304 VDPWR.n158 VDPWR.n157 0.0624718
R1305 VDPWR.n103 VDPWR.n102 0.0612059
R1306 VDPWR.n188 VDPWR 0.0605
R1307 VDPWR.n211 VDPWR 0.0605
R1308 VDPWR VDPWR.n209 0.0605
R1309 VDPWR.n194 VDPWR 0.0605
R1310 VDPWR VDPWR.n181 0.0605
R1311 VDPWR.n104 VDPWR.n103 0.0599468
R1312 VDPWR.n244 VDPWR.n3 0.0577377
R1313 VDPWR.n105 VDPWR.n104 0.0571702
R1314 VDPWR.n106 VDPWR.n105 0.0555
R1315 VDPWR.n107 VDPWR.n106 0.0535722
R1316 VDPWR.n240 VDPWR.n239 0.0532395
R1317 VDPWR.n249 VDPWR.n248 0.0522
R1318 VDPWR.n138 VDPWR.n32 0.0521569
R1319 VDPWR.n108 VDPWR.n107 0.0509772
R1320 VDPWR.n109 VDPWR.n108 0.0493889
R1321 VDPWR.n162 VDPWR.n160 0.0487018
R1322 VDPWR.n110 VDPWR.n109 0.04758
R1323 VDPWR.n238 VDPWR.n8 0.0460752
R1324 VDPWR.n149 VDPWR.n148 0.045577
R1325 VDPWR.n60 VDPWR.n59 0.0448348
R1326 VDPWR.n112 VDPWR.n111 0.0427745
R1327 VDPWR.n242 VDPWR.n241 0.0419028
R1328 VDPWR.n167 VDPWR.n166 0.0415667
R1329 VDPWR.n158 VDPWR.n8 0.0413571
R1330 VDPWR.n244 VDPWR.n243 0.0410333
R1331 VDPWR.n238 VDPWR.n237 0.0408577
R1332 VDPWR.n113 VDPWR.n112 0.0408512
R1333 VDPWR.n183 VDPWR.n174 0.0405
R1334 VDPWR.n155 VDPWR.n9 0.0403491
R1335 VDPWR.n157 VDPWR.n154 0.040162
R1336 VDPWR.n154 VDPWR.n13 0.040162
R1337 VDPWR.n166 VDPWR.n17 0.0397857
R1338 VDPWR.n114 VDPWR.n113 0.0389466
R1339 VDPWR.n166 VDPWR.n165 0.0385976
R1340 VDPWR.n146 VDPWR.n25 0.0383925
R1341 VDPWR.n115 VDPWR.n114 0.0377308
R1342 VDPWR.n148 VDPWR.n25 0.0376329
R1343 VDPWR.n116 VDPWR.n115 0.0358684
R1344 VDPWR.n245 VDPWR.n244 0.0356133
R1345 VDPWR.n237 VDPWR.n9 0.0341226
R1346 VDPWR.n117 VDPWR.n116 0.0338649
R1347 VDPWR.n118 VDPWR.n117 0.0320472
R1348 VDPWR.n119 VDPWR.n118 0.0306596
R1349 VDPWR.n229 VDPWR.n174 0.0305
R1350 VDPWR.n120 VDPWR.n119 0.0288738
R1351 VDPWR.n152 VDPWR.n21 0.0282619
R1352 VDPWR.n121 VDPWR.n120 0.0271047
R1353 VDPWR.n209 VDPWR.n208 0.02675
R1354 VDPWR.n191 VDPWR.n181 0.02675
R1355 VDPWR.n122 VDPWR.n121 0.0257593
R1356 VDPWR.n223 VDPWR.n199 0.0255
R1357 VDPWR.n169 VDPWR.n168 0.0249162
R1358 VDPWR.n235 VDPWR.n11 0.0249162
R1359 VDPWR.n235 VDPWR.n12 0.0249162
R1360 VDPWR.n123 VDPWR.n122 0.0239128
R1361 VDPWR.n136 VDPWR.n135 0.02261
R1362 VDPWR.n124 VDPWR.n123 0.0222982
R1363 VDPWR.n20 VDPWR.n15 0.02162
R1364 VDPWR.n172 VDPWR.n15 0.02162
R1365 VDPWR.n234 VDPWR.n233 0.02162
R1366 VDPWR.n160 VDPWR.n159 0.0212984
R1367 VDPWR.n125 VDPWR.n124 0.0205913
R1368 VDPWR.n126 VDPWR.n125 0.018984
R1369 VDPWR.n241 VDPWR.n4 0.0188236
R1370 VDPWR.n152 VDPWR.n151 0.0182408
R1371 VDPWR.n135 VDPWR.n134 0.0179271
R1372 VDPWR.n127 VDPWR.n126 0.0176222
R1373 VDPWR.n128 VDPWR.n127 0.0160294
R1374 VDPWR.n248 VDPWR.n247 0.015852
R1375 VDPWR.n4 VDPWR.n3 0.0156247
R1376 VDPWR.n240 VDPWR.n6 0.0149236
R1377 VDPWR.n246 VDPWR.n3 0.0148367
R1378 VDPWR.n129 VDPWR.n128 0.0140385
R1379 VDPWR.n156 VDPWR.n14 0.0138871
R1380 VDPWR.n14 VDPWR.n11 0.0133938
R1381 VDPWR.n153 VDPWR.n22 0.0132264
R1382 VDPWR.n171 VDPWR.n16 0.0132264
R1383 VDPWR.n130 VDPWR.n129 0.0131847
R1384 VDPWR.n168 VDPWR.n22 0.0131568
R1385 VDPWR.n169 VDPWR.n16 0.0131568
R1386 VDPWR.n166 VDPWR.n21 0.0115
R1387 VDPWR.n131 VDPWR.n130 0.0112027
R1388 VDPWR.n236 VDPWR.n10 0.0100472
R1389 VDPWR.n13 VDPWR.n10 0.0100023
R1390 VDPWR.n132 VDPWR.n131 0.00957623
R1391 VDPWR.n133 VDPWR.n132 0.00839238
R1392 VDPWR.n237 VDPWR.n236 0.00672642
R1393 VDPWR.n200 VDPWR.n173 0.00661111
R1394 VDPWR.n134 VDPWR.n133 0.00641928
R1395 VDPWR.n159 VDPWR.n10 0.00463323
R1396 VDPWR.n228 VDPWR.n227 0.003
R1397 VDPWR.n197 VDPWR.n195 0.00197617
R1398 VDPWR.n246 VDPWR.n245 0.00108355
R1399 VDPWR.t10 VDPWR.n195 0.00102381
R1400 VDPWR.n202 VDPWR.n198 0.001
R1401 VDPWR.n201 VDPWR.n198 0.001
R1402 VDPWR.t23 VDPWR.n202 0.001
R1403 VDPWR.n201 VDPWR.n197 0.001
R1404 uo_out[2].n3 uo_out[2].t2 15.0005
R1405 uo_out[2] uo_out[2].n3 12.8496
R1406 uo_out[2].n2 uo_out[2] 12.5614
R1407 uo_out[2].n2 uo_out[2].n1 9.01936
R1408 uo_out[2].n0 uo_out[2].t1 8.53421
R1409 uo_out[2].n0 uo_out[2].t0 6.13626
R1410 uo_out[2].n1 uo_out[2].n0 0.0993764
R1411 uo_out[2].n1 uo_out[2] 0.0598258
R1412 uo_out[2] uo_out[2].n2 0.0388429
R1413 uo_out[2].n3 uo_out[2] 0.02525
R1414 uo_out[0].n4 uo_out[0].n3 33.1637
R1415 uo_out[0].n5 uo_out[0].t1 18.0455
R1416 uo_out[0] uo_out[0].t0 18.0125
R1417 uo_out[0].n1 uo_out[0].t3 15.0005
R1418 uo_out[0].n2 uo_out[0].n1 9.03505
R1419 uo_out[0].n3 uo_out[0].n2 6.7505
R1420 uo_out[0].n5 uo_out[0].n4 6.67645
R1421 uo_out[0].n4 uo_out[0].n0 4.90955
R1422 uo_out[0].n0 uo_out[0].t2 3.93974
R1423 uo_out[0].n3 uo_out[0] 1.35863
R1424 uo_out[0] uo_out[0].n5 0.0885
R1425 uo_out[0].n0 uo_out[0] 0.0446962
R1426 uo_out[0].n2 uo_out[0] 0.0401
R1427 uo_out[0].n1 uo_out[0] 0.02525
R1428 uo_out[3].n2 uo_out[3] 15.6957
R1429 uo_out[3].n2 uo_out[3].n1 9.0225
R1430 uo_out[3].n0 uo_out[3].t1 8.53421
R1431 uo_out[3].n0 uo_out[3].t0 6.13626
R1432 uo_out[3].n1 uo_out[3].n0 0.11668
R1433 uo_out[3].n1 uo_out[3] 0.0425225
R1434 uo_out[3] uo_out[3].n2 0.0357
C10 uo_out[0] VGND 11.2531f
C11 VDPWR VGND 0.10244p
.ends

