* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] VAPWR
+ VDPWR VGND
X0 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VAPWR.t25 VAPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X1 VGND.t22 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_5.A VGND.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X2 VDPWR.t51 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_10715_43723# VDPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X3 a_10544_44089# a_10297_43723# VDPWR.t17 VDPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X4 a_10297_43723# a_10168_43997# a_9876_43697# VGND.t77 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X5 a_10368_43697# a_10161_43697# a_10544_44089# VDPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X6 VGND.t48 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X7 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VAPWR.t19 VAPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X8 VGND.t68 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X9 a_13468_43697# a_13740_43697# VGND.t83 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VDPWR.t59 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12647_43723# VDPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X11 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X12 VGND.t1 a_11441_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X13 VAPWR.t9 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VAPWR.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X14 a_12093_43697# uo_out[1].t2 VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X15 a_12051_44089# a_11536_43697# VDPWR.t41 VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X16 VAPWR.t35 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VAPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X17 a_14232_43697# a_14032_43997# a_14381_43723# VGND.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X18 VGND.t11 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X19 VGND.t54 a_13468_43697# uo_out[1].t0 VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X20 VDPWR.t5 a_9509_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X21 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VGND.t82 VGND.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X22 ring_0/skullfet_inverter_9.A skullfet_level_shifter.A VAPWR.t13 VAPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X23 a_13960_43723# a_13468_43697# VGND.t52 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X24 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t85 VGND.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X25 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t87 VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X26 VGND.t95 a_9604_43697# uo_out[3].t0 VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X27 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t89 VGND.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X28 VAPWR.t43 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VAPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X29 VGND.t3 a_14232_43697# a_14161_43723# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X30 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VAPWR.t23 VAPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X31 VGND.t40 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X32 VGND.t5 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X33 a_12647_43723# a_12100_43997# a_12300_43697# VDPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X34 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t46 VGND.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X35 a_13468_43697# a_13740_43697# VDPWR.t61 VDPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X36 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VAPWR.t17 VAPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X37 a_11441_43697# a_11536_43697# VDPWR.t39 VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X38 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t79 VGND.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X39 VDPWR.t48 a_10161_43697# a_10168_43997# VDPWR.t47 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X40 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_5.A VAPWR.t27 VAPWR.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X41 uo_out[0].t0 skullfet_level_shifter.A VGND.t26 VGND.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X42 a_14025_43697# uo_out[0].t2 VGND.t31 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X43 a_14232_43697# a_14025_43697# a_14408_44089# VDPWR.t55 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X44 a_14161_43723# a_14025_43697# a_13740_43697# VDPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X45 VDPWR.t35 a_13468_43697# uo_out[1].t1 VDPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X46 VDPWR.t45 a_12093_43697# a_12100_43997# VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X47 VDPWR.t67 a_9604_43697# uo_out[3].t1 VDPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X48 VGND.t75 a_14025_43697# a_14032_43997# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X49 a_9509_43697# a_9604_43697# VDPWR.t65 VDPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X50 VGND.t9 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X51 a_10119_44089# a_9604_43697# VDPWR.t63 VDPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X52 a_10161_43697# uo_out[2].t2 VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X53 a_13740_43697# a_14032_43997# a_13983_44089# VDPWR.t9 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X54 ua[0].t0 uo_out[0].t3 VAPWR.t31 VAPWR.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X55 VAPWR.t21 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VAPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X56 VGND.t42 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X57 a_12028_43723# a_11536_43697# VGND.t60 VGND.t59 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X58 skullfet_level_shifter.A ring_0/skullfet_inverter_7.A VAPWR.t29 VAPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X59 a_10517_43723# a_10297_43723# VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X60 VAPWR.t41 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VAPWR.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X61 VGND.t70 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_6.A VGND.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X62 a_9604_43697# a_9876_43697# VGND.t37 VGND.t36 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 VGND.t30 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_14579_43723# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X64 a_12093_43697# uo_out[1].t3 VGND.t29 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 VAPWR.t33 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VAPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X66 a_12449_43723# a_12229_43723# VGND.t100 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X67 VGND.t58 a_11536_43697# uo_out[2].t0 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VGND.t7 a_9509_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X69 VGND.t44 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X70 VGND.t38 a_12300_43697# a_12229_43723# VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X71 a_10715_43723# a_10168_43997# a_10368_43697# VDPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X72 a_9604_43697# a_9876_43697# VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X73 a_11536_43697# a_11808_43697# VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X74 a_13373_43697# a_13468_43697# VGND.t51 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X75 a_14408_44089# a_14161_43723# VDPWR.t7 VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X76 VGND.t72 ring_0/skullfet_inverter_7.A skullfet_level_shifter.A VGND.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X77 VGND.t66 a_10161_43697# a_10168_43997# VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X78 a_10096_43723# a_9604_43697# VGND.t93 VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X79 VDPWR.t37 a_11536_43697# uo_out[2].t1 VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X80 VDPWR.t69 a_13373_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X81 VDPWR.t19 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_14579_43723# VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X82 VGND.t62 a_12093_43697# a_12100_43997# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X83 a_14579_43723# a_14025_43697# a_14232_43697# VGND.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X84 a_14161_43723# a_14032_43997# a_13740_43697# VGND.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X85 a_11808_43697# a_12100_43997# a_12051_44089# VDPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X86 VAPWR.t39 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VAPWR.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X87 a_10161_43697# uo_out[2].t3 VGND.t20 VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X88 VAPWR.t37 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VAPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X89 a_10368_43697# a_10168_43997# a_10517_43723# VGND.t76 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X90 a_11536_43697# a_11808_43697# VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X91 VGND.t50 a_10368_43697# a_10297_43723# VGND.t49 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X92 a_12300_43697# a_12100_43997# a_12449_43723# VGND.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X93 a_11808_43697# a_12093_43697# a_12028_43723# VGND.t61 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X94 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VAPWR.t7 VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X95 VDPWR.t13 skullfet_level_shifter.A uo_out[0].t1 VDPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X96 a_13373_43697# a_13468_43697# VDPWR.t33 VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X97 VDPWR.t3 a_14232_43697# a_14161_43723# VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X98 a_13740_43697# a_14025_43697# a_13960_43723# VGND.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X99 a_10297_43723# a_10161_43697# a_9876_43697# VDPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X100 a_11441_43697# a_11536_43697# VGND.t56 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X101 a_12476_44089# a_12229_43723# VDPWR.t73 VDPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X102 a_12229_43723# a_12100_43997# a_11808_43697# VGND.t99 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X103 a_12229_43723# a_12093_43697# a_11808_43697# VDPWR.t43 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X104 a_12300_43697# a_12093_43697# a_12476_44089# VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X105 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VAPWR.t15 VAPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X106 a_10715_43723# a_10161_43697# a_10368_43697# VGND.t64 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X107 VDPWR.t1 a_11441_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X108 VGND.t15 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X109 VGND.t24 skullfet_level_shifter.A ring_0/skullfet_inverter_9.A VGND.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X110 VGND.t98 a_13373_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X111 a_9509_43697# a_9604_43697# VGND.t91 VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X112 VGND.t74 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_10715_43723# VGND.t73 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X113 a_12647_43723# a_12093_43697# a_12300_43697# VGND.t16 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X114 a_9876_43697# a_10168_43997# a_10119_44089# VDPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X115 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_4.A VAPWR.t11 VAPWR.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X116 a_14381_43723# a_14161_43723# VGND.t13 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X117 VGND.t80 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12647_43723# VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X118 VGND.t35 uo_out[0].t4 ua[0].t1 VGND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X119 a_14579_43723# a_14032_43997# a_14232_43697# VDPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X120 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VGND.t18 VGND.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X121 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VAPWR.t3 VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X122 VDPWR.t29 a_10368_43697# a_10297_43723# VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X123 a_9876_43697# a_10161_43697# a_10096_43723# VGND.t63 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X124 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VAPWR.t5 VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X125 a_14025_43697# uo_out[0].t5 VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X126 a_13983_44089# a_13468_43697# VDPWR.t31 VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X127 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t97 VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X128 VDPWR.t27 a_12300_43697# a_12229_43723# VDPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X129 VDPWR.t53 a_14025_43697# a_14032_43997# VDPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
R0 VAPWR.n68 VAPWR.t31 738.801
R1 VAPWR.n52 VAPWR.t21 738.799
R2 VAPWR.n54 VAPWR.t23 738.799
R3 VAPWR.n38 VAPWR.t9 738.799
R4 VAPWR.n34 VAPWR.t35 738.799
R5 VAPWR.n6 VAPWR.t17 738.799
R6 VAPWR.n41 VAPWR.t41 738.799
R7 VAPWR.n44 VAPWR.t39 738.799
R8 VAPWR.n47 VAPWR.t37 738.799
R9 VAPWR.n4 VAPWR.t33 738.799
R10 VAPWR.n2 VAPWR.t43 738.799
R11 VAPWR.n60 VAPWR.t3 738.799
R12 VAPWR.n57 VAPWR.t15 738.799
R13 VAPWR.n32 VAPWR.t7 738.799
R14 VAPWR.n7 VAPWR.t1 738.799
R15 VAPWR.n11 VAPWR.t27 738.799
R16 VAPWR.n22 VAPWR.t25 738.799
R17 VAPWR.n19 VAPWR.t29 738.799
R18 VAPWR.n16 VAPWR.t13 738.799
R19 VAPWR.n13 VAPWR.t5 738.799
R20 VAPWR.n9 VAPWR.t11 738.799
R21 VAPWR.n27 VAPWR.t19 738.799
R22 VAPWR.n68 VAPWR.t30 707.519
R23 VAPWR.n60 VAPWR.t2 707.519
R24 VAPWR.n57 VAPWR.t14 707.519
R25 VAPWR.n52 VAPWR.t20 707.519
R26 VAPWR.n54 VAPWR.t22 707.519
R27 VAPWR.n38 VAPWR.t8 707.519
R28 VAPWR.n34 VAPWR.t34 707.519
R29 VAPWR.n32 VAPWR.t6 707.519
R30 VAPWR.n6 VAPWR.t16 707.519
R31 VAPWR.n7 VAPWR.t0 707.519
R32 VAPWR.n11 VAPWR.t26 707.519
R33 VAPWR.n22 VAPWR.t24 707.519
R34 VAPWR.n19 VAPWR.t28 707.519
R35 VAPWR.n16 VAPWR.t12 707.519
R36 VAPWR.n13 VAPWR.t4 707.519
R37 VAPWR.n9 VAPWR.t10 707.519
R38 VAPWR.n27 VAPWR.t18 707.519
R39 VAPWR.n41 VAPWR.t40 707.519
R40 VAPWR.n44 VAPWR.t38 707.519
R41 VAPWR.n47 VAPWR.t36 707.519
R42 VAPWR.n4 VAPWR.t32 707.519
R43 VAPWR.n2 VAPWR.t42 707.519
R44 VAPWR.n69 VAPWR.n68 13.3797
R45 VAPWR.n61 VAPWR.n60 13.3797
R46 VAPWR.n58 VAPWR.n57 13.3797
R47 VAPWR.n33 VAPWR.n32 13.3797
R48 VAPWR.n8 VAPWR.n7 13.3797
R49 VAPWR.n12 VAPWR.n11 13.3797
R50 VAPWR.n23 VAPWR.n22 13.3797
R51 VAPWR.n20 VAPWR.n19 13.3797
R52 VAPWR.n17 VAPWR.n16 13.3797
R53 VAPWR.n14 VAPWR.n13 13.3797
R54 VAPWR.n10 VAPWR.n9 13.3797
R55 VAPWR.n28 VAPWR.n27 13.3797
R56 VAPWR.n53 VAPWR.n52 13.3223
R57 VAPWR VAPWR.n54 13.3223
R58 VAPWR.n39 VAPWR.n38 13.3223
R59 VAPWR.n35 VAPWR.n34 13.3223
R60 VAPWR VAPWR.n6 13.3223
R61 VAPWR.n42 VAPWR.n41 13.3223
R62 VAPWR.n45 VAPWR.n44 13.3223
R63 VAPWR.n48 VAPWR.n47 13.3223
R64 VAPWR.n5 VAPWR.n4 13.3223
R65 VAPWR.n3 VAPWR.n2 13.3223
R66 VAPWR.n70 VAPWR.n69 10.0371
R67 VAPWR.n59 VAPWR.n58 9.70762
R68 VAPWR.n18 VAPWR.n15 9.45042
R69 VAPWR.n31 VAPWR 8.52916
R70 VAPWR.n62 VAPWR.n61 7.92611
R71 VAPWR.n40 VAPWR.n37 7.71912
R72 VAPWR.n15 VAPWR.n14 7.71771
R73 VAPWR.n31 VAPWR.n30 7.41572
R74 VAPWR.n55 VAPWR 7.13154
R75 VAPWR.n40 VAPWR.n39 7.11663
R76 VAPWR.n18 VAPWR.n17 7.10884
R77 VAPWR.n43 VAPWR.n42 6.89753
R78 VAPWR.n21 VAPWR.n20 6.54898
R79 VAPWR.n49 VAPWR.n46 6.23852
R80 VAPWR.n30 VAPWR.n8 6.19396
R81 VAPWR.n46 VAPWR.n45 6.10554
R82 VAPWR.n29 VAPWR.n28 6.01845
R83 VAPWR.n36 VAPWR.n35 5.92055
R84 VAPWR.n49 VAPWR.n48 5.84717
R85 VAPWR.n24 VAPWR.n23 5.78073
R86 VAPWR.n26 VAPWR.n10 5.73072
R87 VAPWR.n50 VAPWR.n5 5.60146
R88 VAPWR.n51 VAPWR.n3 5.59565
R89 VAPWR.n25 VAPWR.n12 5.50466
R90 VAPWR.n55 VAPWR.n53 4.89777
R91 VAPWR.n36 VAPWR.n33 4.86074
R92 VAPWR.n46 VAPWR.n43 4.01511
R93 VAPWR.n66 VAPWR 3.49767
R94 VAPWR.n70 VAPWR.n67 3.40236
R95 VAPWR.n37 VAPWR.n36 2.91269
R96 VAPWR.n59 VAPWR.n56 2.82184
R97 VAPWR.n1 VAPWR.n0 1.63622
R98 VAPWR.n24 VAPWR.n21 1.36014
R99 VAPWR.n30 VAPWR.n29 1.34127
R100 VAPWR.n56 VAPWR.n51 1.32921
R101 VAPWR.n56 VAPWR.n55 1.313
R102 VAPWR.n63 VAPWR.n0 1.29727
R103 VAPWR.n29 VAPWR.n26 1.10191
R104 VAPWR.n51 VAPWR.n50 0.940035
R105 VAPWR.n62 VAPWR.n59 0.85748
R106 VAPWR.n37 VAPWR.n31 0.767594
R107 VAPWR.n66 VAPWR.n65 0.616014
R108 VAPWR.n25 VAPWR.n24 0.52495
R109 VAPWR.n43 VAPWR.n40 0.514977
R110 VAPWR.n15 VAPWR.n1 0.507476
R111 VAPWR.n26 VAPWR.n25 0.505442
R112 VAPWR.n21 VAPWR.n18 0.500622
R113 VAPWR.n50 VAPWR.n49 0.483622
R114 VAPWR.n65 VAPWR.n0 0.20333
R115 VAPWR.n67 VAPWR 0.193138
R116 VAPWR.n69 VAPWR 0.057877
R117 VAPWR.n61 VAPWR 0.057877
R118 VAPWR.n58 VAPWR 0.057877
R119 VAPWR.n33 VAPWR 0.057877
R120 VAPWR.n8 VAPWR 0.057877
R121 VAPWR.n12 VAPWR 0.057877
R122 VAPWR.n23 VAPWR 0.057877
R123 VAPWR.n20 VAPWR 0.057877
R124 VAPWR.n17 VAPWR 0.057877
R125 VAPWR.n14 VAPWR 0.057877
R126 VAPWR.n10 VAPWR 0.057877
R127 VAPWR.n28 VAPWR 0.057877
R128 VAPWR.n53 VAPWR 0.0496071
R129 VAPWR.n39 VAPWR 0.0496071
R130 VAPWR.n35 VAPWR 0.0496071
R131 VAPWR.n42 VAPWR 0.0496071
R132 VAPWR.n45 VAPWR 0.0496071
R133 VAPWR.n48 VAPWR 0.0496071
R134 VAPWR.n5 VAPWR 0.0496071
R135 VAPWR.n3 VAPWR 0.0496071
R136 VAPWR VAPWR.n70 0.0475
R137 VAPWR.n65 VAPWR.n64 0.0335189
R138 VAPWR.n70 VAPWR 0.024
R139 VAPWR.n64 VAPWR.n1 0.00474612
R140 VAPWR.n63 VAPWR.n62 0.00305102
R141 VAPWR.n64 VAPWR.n63 0.00285849
R142 VAPWR.n67 VAPWR.n66 0.0018126
R143 VGND.n394 VGND.n393 101372
R144 VGND.n408 VGND.n407 97829.8
R145 VGND.n452 VGND.n10 64989.2
R146 VGND.n392 VGND.n391 63317.7
R147 VGND.n320 VGND.n315 49981.2
R148 VGND.n329 VGND.t8 48989.1
R149 VGND.n390 VGND.n317 48956.8
R150 VGND.n236 VGND.n15 46397.1
R151 VGND.n318 VGND.n29 34056.2
R152 VGND.t67 VGND.n27 32820.9
R153 VGND.n355 VGND.n352 31013.9
R154 VGND.n358 VGND.n352 30664.6
R155 VGND.n143 VGND.n27 30664.6
R156 VGND.n410 VGND.n409 29705.2
R157 VGND.n321 VGND.n320 26125.9
R158 VGND.n330 VGND.n329 24501.8
R159 VGND.n332 VGND.n321 22668.4
R160 VGND.n393 VGND.n317 20954.6
R161 VGND.n407 VGND.n29 20954.6
R162 VGND.n409 VGND.n408 20954.6
R163 VGND.n323 VGND.n13 18294.4
R164 VGND.t6 VGND.n15 14642.2
R165 VGND.n352 VGND.n317 13862.9
R166 VGND.n409 VGND.n27 13853.3
R167 VGND.n312 VGND.n310 13669.6
R168 VGND.n329 VGND.n321 10983.3
R169 VGND.n236 VGND.n235 10461.7
R170 VGND.n391 VGND.t45 8761.83
R171 VGND.n332 VGND.n331 8254.98
R172 VGND.n408 VGND.n10 8171.07
R173 VGND.n393 VGND.n392 8164.43
R174 VGND.n453 VGND.n452 8158.04
R175 VGND.n452 VGND.n13 8007.21
R176 VGND.n391 VGND.n332 8000.6
R177 VGND.n406 VGND.n31 7798.05
R178 VGND.n236 VGND 7183.82
R179 VGND.n310 VGND.n31 7076.09
R180 VGND.n392 VGND.n320 6658.85
R181 VGND.n13 VGND.n12 6298.11
R182 VGND.n391 VGND.n390 5608.83
R183 VGND.n238 VGND.n237 5446.6
R184 VGND.n312 VGND.n311 4952.1
R185 VGND.n318 VGND.n10 4690.48
R186 VGND.n400 VGND.t14 4526.67
R187 VGND.n395 VGND.n315 4456.64
R188 VGND.n330 VGND.n322 4323.23
R189 VGND.n326 VGND.n13 4311.21
R190 VGND.n405 VGND.t14 3320.6
R191 VGND.n319 VGND.n31 3097.77
R192 VGND.n323 VGND.n320 3097.77
R193 VGND.n396 VGND.n314 3043.22
R194 VGND.n326 VGND.n325 2374.28
R195 VGND.n328 VGND.n326 2325.64
R196 VGND.n394 VGND.t88 2293.69
R197 VGND.n452 VGND.n14 2139.51
R198 VGND.n384 VGND.t45 2108.34
R199 VGND.n396 VGND.n31 2021.45
R200 VGND.t17 VGND.n314 1523.34
R201 VGND.n12 VGND.t10 1523.34
R202 VGND.n453 VGND.t23 1523.34
R203 VGND.n407 VGND.t43 1467.82
R204 VGND.n406 VGND.n30 1463.87
R205 VGND.n390 VGND.t96 1206.01
R206 VGND.n414 VGND.n413 1198.25
R207 VGND.n412 VGND.n25 1198.25
R208 VGND.n311 VGND.n0 963.163
R209 VGND.n306 VGND.n29 921.593
R210 VGND.n359 VGND.n316 892.495
R211 VGND.n389 VGND.t78 842.21
R212 VGND.t92 VGND.t36 809.293
R213 VGND.n407 VGND.n406 807.846
R214 VGND.t94 VGND.t90 800.774
R215 VGND.t21 VGND.n28 787.793
R216 VGND.n310 VGND.t14 759.1
R217 VGND.n395 VGND.n394 634.295
R218 VGND.n311 VGND.t34 614.494
R219 VGND.n451 VGND.n15 613.852
R220 VGND.n235 VGND.n234 595.942
R221 VGND.n30 VGND.n29 587.612
R222 VGND.n314 VGND.n313 585
R223 VGND.n12 VGND.n11 585
R224 VGND.n328 VGND.n327 585
R225 VGND.n451 VGND.n450 585
R226 VGND.n357 VGND.n356 585
R227 VGND.n354 VGND.n353 585
R228 VGND.n389 VGND.n388 585
R229 VGND.n361 VGND.n316 585
R230 VGND.n360 VGND.n359 585
R231 VGND.n398 VGND.n397 585
R232 VGND.n325 VGND.n324 585
R233 VGND.n454 VGND.n453 585
R234 VGND.n74 VGND.n14 585
R235 VGND.n146 VGND.n145 585
R236 VGND.n239 VGND.n238 585
R237 VGND.n33 VGND.n28 585
R238 VGND.n142 VGND.n141 585
R239 VGND.n405 VGND.n404 585
R240 VGND.t8 VGND.n328 574.539
R241 VGND.t69 VGND.n143 539.317
R242 VGND.t84 VGND.n355 533.332
R243 VGND.t86 VGND.n358 500.077
R244 VGND.n238 VGND.t67 489.839
R245 VGND.t77 VGND.t63 451.5
R246 VGND.t49 VGND.t77 430.204
R247 VGND.n30 VGND.t4 427.527
R248 VGND.n331 VGND.t47 424.175
R249 VGND.t63 VGND.t92 404.647
R250 VGND.t90 VGND.t6 404.647
R251 VGND.n355 VGND.n354 382.728
R252 VGND.n143 VGND.n142 377.945
R253 VGND.n411 VGND.t49 370.572
R254 VGND.n325 VGND.t39 362.452
R255 VGND.n315 VGND.t17 360.884
R256 VGND.n358 VGND.n357 360.842
R257 VGND.t36 VGND.t94 357.793
R258 VGND.n452 VGND.t25 313.435
R259 VGND.n407 VGND.n28 302.216
R260 VGND.n0 VGND.t35 282.132
R261 VGND.n239 VGND.t68 282.13
R262 VGND.n306 VGND.t5 282.13
R263 VGND.n141 VGND.t22 282.13
R264 VGND.n33 VGND.t44 282.13
R265 VGND.n11 VGND.t11 282.13
R266 VGND.n327 VGND.t9 282.13
R267 VGND.n400 VGND.t15 282.13
R268 VGND.n324 VGND.t40 282.13
R269 VGND.n454 VGND.t24 282.13
R270 VGND.n74 VGND.t72 282.13
R271 VGND.n145 VGND.t70 282.13
R272 VGND.n450 VGND.t26 281.841
R273 VGND.n404 VGND.t42 281.839
R274 VGND.n398 VGND.t82 281.839
R275 VGND.n360 VGND.t87 281.839
R276 VGND.n361 VGND.t89 281.839
R277 VGND.n384 VGND.t46 281.839
R278 VGND.n313 VGND.t18 281.839
R279 VGND.n322 VGND.t48 281.839
R280 VGND.n388 VGND.t97 281.839
R281 VGND.n353 VGND.t79 281.839
R282 VGND.n356 VGND.t85 281.839
R283 VGND.n329 VGND.n323 264.286
R284 VGND.n177 VGND.t52 251
R285 VGND.n214 VGND.t60 251
R286 VGND.n437 VGND.t93 251
R287 VGND.n331 VGND.t39 245.631
R288 VGND.n157 VGND.t30 243.028
R289 VGND.n227 VGND.t80 243.028
R290 VGND.n424 VGND.t74 243.028
R291 VGND.n411 VGND.t71 232.994
R292 VGND.n179 VGND.n151 218.506
R293 VGND.n201 VGND.n200 218.506
R294 VGND.n439 VGND.n438 218.506
R295 VGND.t25 VGND.n451 212.357
R296 VGND.n320 VGND.n319 209.014
R297 VGND.n186 VGND.n185 200.201
R298 VGND.n204 VGND.n203 200.201
R299 VGND.n447 VGND.n446 200.201
R300 VGND.n160 VGND.n159 199.739
R301 VGND.n192 VGND.n191 199.739
R302 VGND.n420 VGND.n419 199.739
R303 VGND.n155 VGND.n154 199.53
R304 VGND.n221 VGND.n196 199.53
R305 VGND.n430 VGND.n22 199.53
R306 VGND.t71 VGND.n14 196.702
R307 VGND.n396 VGND.n395 178.196
R308 VGND.n237 VGND.n236 165.179
R309 VGND.n146 VGND.t69 162.868
R310 VGND.n142 VGND.t21 153.912
R311 VGND.n357 VGND.t84 153.888
R312 VGND.n354 VGND.t78 151.095
R313 VGND.t96 VGND.n389 151.095
R314 VGND.n359 VGND.t86 145.869
R315 VGND.t81 VGND.n396 130.082
R316 VGND.n406 VGND.t41 129.425
R317 VGND.t16 VGND 118.189
R318 VGND.n397 VGND.t81 99.8351
R319 VGND.t41 VGND.n405 99.332
R320 VGND.n154 VGND.t3 74.8666
R321 VGND.n196 VGND.t38 74.8666
R322 VGND.n22 VGND.t50 74.8666
R323 VGND.n394 VGND.n316 73.7658
R324 VGND.t59 VGND.t32 69.615
R325 VGND.t57 VGND.t55 68.8822
R326 VGND.t65 VGND.t73 68.8822
R327 VGND.t47 VGND.n330 54.4208
R328 VGND.n185 VGND.t51 54.2862
R329 VGND.n203 VGND.t56 54.2862
R330 VGND.n446 VGND.t91 54.2862
R331 VGND.n397 VGND.n312 54.1077
R332 VGND.n236 VGND.n146 53.7948
R333 VGND.t73 VGND.t64 41.0364
R334 VGND.n154 VGND.t13 40.0005
R335 VGND.n196 VGND.t100 40.0005
R336 VGND.n22 VGND.t28 40.0005
R337 VGND.t99 VGND.t61 38.838
R338 VGND.n159 VGND.t31 38.5719
R339 VGND.n159 VGND.t75 38.5719
R340 VGND.n191 VGND.t29 38.5719
R341 VGND.n191 VGND.t62 38.5719
R342 VGND.n419 VGND.t20 38.5719
R343 VGND.n419 VGND.t66 38.5719
R344 VGND.t64 VGND.t76 36.2733
R345 VGND.t76 VGND.t27 36.2733
R346 VGND.t61 VGND.t59 34.8077
R347 VGND.t55 VGND.t0 34.8077
R348 VGND.n166 VGND.n165 34.6358
R349 VGND.n167 VGND.n166 34.6358
R350 VGND.n172 VGND.n171 34.6358
R351 VGND.n173 VGND.n172 34.6358
R352 VGND.n173 VGND.n152 34.6358
R353 VGND.n180 VGND.n149 34.6358
R354 VGND.n184 VGND.n149 34.6358
R355 VGND.n226 VGND.n194 34.6358
R356 VGND.n222 VGND.n194 34.6358
R357 VGND.n220 VGND.n197 34.6358
R358 VGND.n216 VGND.n197 34.6358
R359 VGND.n216 VGND.n215 34.6358
R360 VGND.n210 VGND.n209 34.6358
R361 VGND.n209 VGND.n208 34.6358
R362 VGND.n426 VGND.n425 34.6358
R363 VGND.n426 VGND.n21 34.6358
R364 VGND.n432 VGND.n431 34.6358
R365 VGND.n432 VGND.n19 34.6358
R366 VGND.n436 VGND.n19 34.6358
R367 VGND.n444 VGND.n17 34.6358
R368 VGND.n445 VGND.n444 34.6358
R369 VGND.n413 VGND.n412 33.7085
R370 VGND.n412 VGND 33.7085
R371 VGND.n179 VGND.n178 32.7534
R372 VGND.n213 VGND.n201 32.7534
R373 VGND.n440 VGND.n439 32.7534
R374 VGND.t2 VGND.t12 31.3274
R375 VGND.n178 VGND.n177 31.2476
R376 VGND.n214 VGND.n213 31.2476
R377 VGND.n440 VGND.n437 31.2476
R378 VGND.n167 VGND.n155 30.8711
R379 VGND.n222 VGND.n221 30.8711
R380 VGND.n430 VGND.n21 30.8711
R381 VGND.t32 VGND.t57 30.7774
R382 VGND.t19 VGND.t65 30.7774
R383 VGND.n165 VGND.n157 27.4829
R384 VGND.n227 VGND.n226 27.4829
R385 VGND.n425 VGND.n424 27.4829
R386 VGND.n185 VGND.t98 25.9346
R387 VGND.n203 VGND.t1 25.9346
R388 VGND.n446 VGND.t7 25.9346
R389 VGND.n410 VGND.t0 25.6479
R390 VGND.n413 VGND.n410 25.6479
R391 VGND.n151 VGND.t83 24.9236
R392 VGND.n151 VGND.t54 24.9236
R393 VGND.n200 VGND.t33 24.9236
R394 VGND.n200 VGND.t58 24.9236
R395 VGND.n438 VGND.t37 24.9236
R396 VGND.n438 VGND.t95 24.9236
R397 VGND.n362 VGND.n309 23.8781
R398 VGND.n186 VGND.n184 23.7181
R399 VGND.n187 VGND.n147 23.7181
R400 VGND.n233 VGND.n232 23.7181
R401 VGND.n208 VGND.n204 23.7181
R402 VGND.n414 VGND.n26 23.7181
R403 VGND.n418 VGND.n25 23.7181
R404 VGND.n447 VGND.n445 23.7181
R405 VGND.n385 VGND.n2 23.1263
R406 VGND.n161 VGND.n160 22.9652
R407 VGND.n161 VGND.n157 22.9652
R408 VGND.n228 VGND.n192 22.9652
R409 VGND.n228 VGND.n227 22.9652
R410 VGND.n420 VGND.n24 22.9652
R411 VGND.n424 VGND.n24 22.9652
R412 VGND.n235 VGND.t53 22.7837
R413 VGND.n177 VGND.n152 22.2123
R414 VGND.n215 VGND.n214 22.2123
R415 VGND.n437 VGND.n436 22.2123
R416 VGND.n187 VGND.n186 21.4593
R417 VGND.n232 VGND.n192 21.4593
R418 VGND.n204 VGND.n26 21.4593
R419 VGND.n420 VGND.n418 21.4593
R420 VGND.n462 VGND.n461 20.8917
R421 VGND.n403 VGND.n308 19.445
R422 VGND.n319 VGND.n318 15.7795
R423 VGND.n240 VGND.n239 13.2958
R424 VGND.n307 VGND.n306 13.2958
R425 VGND.n141 VGND.n140 13.2958
R426 VGND.n34 VGND.n33 13.2958
R427 VGND.n11 VGND.n5 13.2958
R428 VGND.n327 VGND.n4 13.2958
R429 VGND.n401 VGND.n400 13.2958
R430 VGND.n324 VGND.n3 13.2958
R431 VGND.n455 VGND.n454 13.2958
R432 VGND.n75 VGND.n74 13.2958
R433 VGND.n145 VGND.n144 13.2958
R434 VGND.n468 VGND.n0 13.2958
R435 VGND.n404 VGND 13.2396
R436 VGND VGND.n398 13.2396
R437 VGND VGND.n361 13.2396
R438 VGND.n313 VGND 13.2396
R439 VGND.n322 VGND 13.2396
R440 VGND.n450 VGND 13.2396
R441 VGND.n388 VGND 13.2396
R442 VGND.n353 VGND 13.2396
R443 VGND.n356 VGND 13.2396
R444 VGND VGND.n384 13.2396
R445 VGND VGND.n360 13.2396
R446 VGND.n237 VGND.t99 13.1906
R447 VGND.n468 VGND 13.1357
R448 VGND VGND.n449 12.8296
R449 VGND.n414 VGND.n25 12.8005
R450 VGND.n449 VGND 12.1807
R451 VGND.t27 VGND.n411 11.725
R452 VGND.n399 VGND.n309 11.3687
R453 VGND VGND.t19 11.3586
R454 VGND.n171 VGND.n155 10.5417
R455 VGND.n221 VGND.n220 10.5417
R456 VGND.n431 VGND.n430 10.5417
R457 VGND.n445 VGND.n16 9.3005
R458 VGND.n444 VGND.n443 9.3005
R459 VGND.n442 VGND.n17 9.3005
R460 VGND.n441 VGND.n440 9.3005
R461 VGND.n437 VGND.n18 9.3005
R462 VGND.n436 VGND.n435 9.3005
R463 VGND.n434 VGND.n19 9.3005
R464 VGND.n433 VGND.n432 9.3005
R465 VGND.n431 VGND.n20 9.3005
R466 VGND.n430 VGND.n429 9.3005
R467 VGND.n428 VGND.n21 9.3005
R468 VGND.n427 VGND.n426 9.3005
R469 VGND.n425 VGND.n23 9.3005
R470 VGND.n424 VGND.n423 9.3005
R471 VGND.n422 VGND.n24 9.3005
R472 VGND.n421 VGND.n420 9.3005
R473 VGND.n418 VGND.n417 9.3005
R474 VGND.n416 VGND.n25 9.3005
R475 VGND.n162 VGND.n161 9.3005
R476 VGND.n163 VGND.n157 9.3005
R477 VGND.n165 VGND.n164 9.3005
R478 VGND.n166 VGND.n156 9.3005
R479 VGND.n168 VGND.n167 9.3005
R480 VGND.n169 VGND.n155 9.3005
R481 VGND.n171 VGND.n170 9.3005
R482 VGND.n172 VGND.n153 9.3005
R483 VGND.n174 VGND.n173 9.3005
R484 VGND.n175 VGND.n152 9.3005
R485 VGND.n177 VGND.n176 9.3005
R486 VGND.n178 VGND.n150 9.3005
R487 VGND.n181 VGND.n180 9.3005
R488 VGND.n182 VGND.n149 9.3005
R489 VGND.n184 VGND.n183 9.3005
R490 VGND.n186 VGND.n148 9.3005
R491 VGND.n188 VGND.n187 9.3005
R492 VGND.n189 VGND.n147 9.3005
R493 VGND.n233 VGND.n190 9.3005
R494 VGND.n232 VGND.n231 9.3005
R495 VGND.n230 VGND.n192 9.3005
R496 VGND.n229 VGND.n228 9.3005
R497 VGND.n227 VGND.n193 9.3005
R498 VGND.n226 VGND.n225 9.3005
R499 VGND.n224 VGND.n194 9.3005
R500 VGND.n223 VGND.n222 9.3005
R501 VGND.n221 VGND.n195 9.3005
R502 VGND.n220 VGND.n219 9.3005
R503 VGND.n218 VGND.n197 9.3005
R504 VGND.n217 VGND.n216 9.3005
R505 VGND.n215 VGND.n198 9.3005
R506 VGND.n214 VGND.n199 9.3005
R507 VGND.n213 VGND.n212 9.3005
R508 VGND.n211 VGND.n210 9.3005
R509 VGND.n209 VGND.n202 9.3005
R510 VGND.n208 VGND.n207 9.3005
R511 VGND.n206 VGND.n204 9.3005
R512 VGND.n205 VGND.n26 9.3005
R513 VGND.n415 VGND.n414 9.3005
R514 VGND VGND.n2 9.06372
R515 VGND.t12 VGND.t16 8.54419
R516 VGND.n402 VGND.n401 7.80496
R517 VGND.n308 VGND.n307 7.42221
R518 VGND.n160 VGND.n158 7.12576
R519 VGND.n448 VGND.n447 7.12063
R520 VGND.n463 VGND.n4 6.96
R521 VGND.n385 VGND 6.82321
R522 VGND.n234 VGND.n147 6.367
R523 VGND.n234 VGND.n233 6.367
R524 VGND.n464 VGND.n3 6.32363
R525 VGND.n304 VGND.n34 6.24462
R526 VGND VGND.n387 6.10287
R527 VGND VGND.n403 5.99098
R528 VGND VGND.n309 5.98182
R529 VGND.n462 VGND.n5 5.94997
R530 VGND.n456 VGND.n455 5.91022
R531 VGND.n362 VGND 5.81859
R532 VGND.n144 VGND.n53 5.80858
R533 VGND.n140 VGND.n43 5.70662
R534 VGND VGND.n351 5.69376
R535 VGND.n363 VGND 5.57954
R536 VGND.n364 VGND 5.53239
R537 VGND.n399 VGND 5.49935
R538 VGND.n121 VGND.n75 5.39911
R539 VGND.n248 VGND.n247 5.04217
R540 VGND.n241 VGND.n240 5.00883
R541 VGND.n449 VGND.n1 4.99159
R542 VGND.n1 VGND 3.44325
R543 VGND VGND.n467 3.36335
R544 VGND.n247 VGND.n246 3.29217
R545 VGND.n308 VGND.n305 3.10947
R546 VGND.n467 VGND 2.3855
R547 VGND.n180 VGND.n179 1.88285
R548 VGND.n210 VGND.n201 1.88285
R549 VGND.n439 VGND.n17 1.88285
R550 VGND.n111 VGND.n110 1.5618
R551 VGND.t53 VGND.t2 1.42445
R552 VGND.n402 VGND.n399 1.28527
R553 VGND.n242 VGND.n241 1.2755
R554 VGND.n249 VGND.n53 0.979021
R555 VGND.n386 VGND.n385 0.96878
R556 VGND.n464 VGND.n463 0.964749
R557 VGND.n403 VGND.n402 0.93288
R558 VGND.n463 VGND.n462 0.903134
R559 VGND.n364 VGND.n363 0.844578
R560 VGND.n110 VGND.n109 0.777168
R561 VGND.n466 VGND.n465 0.726602
R562 VGND.n363 VGND.n362 0.707232
R563 VGND.n247 VGND.n53 0.6755
R564 VGND.n241 VGND.n55 0.638
R565 VGND.n365 VGND.n364 0.577069
R566 VGND.n250 VGND.n249 0.574766
R567 VGND.n465 VGND.n2 0.561048
R568 VGND.n109 VGND.n108 0.533644
R569 VGND.n251 VGND.n250 0.469554
R570 VGND.n251 VGND.n51 0.431514
R571 VGND.n246 VGND.n245 0.425271
R572 VGND.n108 VGND.n107 0.420347
R573 VGND.n107 VGND.n106 0.36938
R574 VGND.n255 VGND.n51 0.355217
R575 VGND.n106 VGND.n105 0.332442
R576 VGND.n256 VGND.n255 0.314827
R577 VGND.n366 VGND.n365 0.307815
R578 VGND.n105 VGND.n104 0.293921
R579 VGND.n257 VGND.n256 0.283145
R580 VGND.n104 VGND.n103 0.262603
R581 VGND.n257 VGND.n49 0.257575
R582 VGND.n103 VGND.n102 0.242676
R583 VGND.n261 VGND.n49 0.242107
R584 VGND.n102 VGND.n101 0.227688
R585 VGND.n262 VGND.n261 0.224203
R586 VGND.n278 VGND.n43 0.21925
R587 VGND.n101 VGND.n100 0.214493
R588 VGND.n263 VGND.n262 0.209128
R589 VGND.n386 VGND.n383 0.207265
R590 VGND.n100 VGND.n96 0.207112
R591 VGND.n101 VGND.n95 0.205418
R592 VGND.n102 VGND.n94 0.203752
R593 VGND.n367 VGND.n366 0.202174
R594 VGND.n100 VGND.n99 0.201991
R595 VGND.n103 VGND.n93 0.2005
R596 VGND.n104 VGND.n92 0.198913
R597 VGND.n105 VGND.n91 0.19735
R598 VGND.n263 VGND.n47 0.196195
R599 VGND.n106 VGND.n90 0.195812
R600 VGND.n99 VGND.n9 0.194723
R601 VGND.n107 VGND.n89 0.194298
R602 VGND.n456 VGND.n8 0.193682
R603 VGND.n108 VGND.n88 0.19134
R604 VGND.n368 VGND.n367 0.190823
R605 VGND.n109 VGND.n87 0.189894
R606 VGND.n267 VGND.n47 0.189066
R607 VGND.n110 VGND.n86 0.18847
R608 VGND.n461 VGND.n6 0.188059
R609 VGND.n369 VGND.n368 0.184664
R610 VGND.n460 VGND.n459 0.181056
R611 VGND.n370 VGND.n369 0.180457
R612 VGND.n268 VGND.n267 0.179109
R613 VGND.n269 VGND.n268 0.178762
R614 VGND.n371 VGND.n370 0.167949
R615 VGND.n269 VGND.n45 0.166149
R616 VGND.n305 VGND.n304 0.165057
R617 VGND.n373 VGND.n372 0.164532
R618 VGND.n372 VGND.n371 0.164276
R619 VGND.n274 VGND.n273 0.159573
R620 VGND.n273 VGND.n45 0.159247
R621 VGND.n139 VGND.n138 0.159247
R622 VGND.n120 VGND.n119 0.156646
R623 VGND.n138 VGND.n137 0.156448
R624 VGND.n374 VGND.n373 0.155102
R625 VGND.n250 VGND.n52 0.154588
R626 VGND.n99 VGND.n98 0.153861
R627 VGND.n252 VGND.n251 0.153802
R628 VGND.n275 VGND.n274 0.153257
R629 VGND.n375 VGND.n374 0.153062
R630 VGND.n253 VGND.n51 0.153016
R631 VGND VGND.n448 0.152603
R632 VGND.n242 VGND.n139 0.152527
R633 VGND.n256 VGND.n50 0.152399
R634 VGND.n245 VGND.n55 0.152332
R635 VGND.n255 VGND.n254 0.15223
R636 VGND.n136 VGND.n135 0.151068
R637 VGND.n259 VGND.n49 0.150816
R638 VGND.n376 VGND.n375 0.150802
R639 VGND.n258 VGND.n257 0.150657
R640 VGND.n137 VGND.n136 0.15035
R641 VGND.n262 VGND.n48 0.150182
R642 VGND.n382 VGND.n334 0.150148
R643 VGND.n261 VGND.n260 0.150025
R644 VGND.n366 VGND.n350 0.149538
R645 VGND.n264 VGND.n263 0.149385
R646 VGND.n368 VGND.n348 0.148887
R647 VGND.n367 VGND.n349 0.148737
R648 VGND.n265 VGND.n47 0.148589
R649 VGND.n448 VGND.n16 0.148519
R650 VGND.n369 VGND.n347 0.148081
R651 VGND.n268 VGND.n46 0.147936
R652 VGND.n267 VGND.n266 0.147793
R653 VGND.n372 VGND.n344 0.147559
R654 VGND.n248 VGND.n54 0.147513
R655 VGND.n371 VGND.n345 0.147416
R656 VGND.n271 VGND.n45 0.147274
R657 VGND.n370 VGND.n346 0.147274
R658 VGND.n139 VGND.n56 0.147274
R659 VGND.n270 VGND.n269 0.147135
R660 VGND.n244 VGND.n243 0.147135
R661 VGND.n375 VGND.n341 0.147023
R662 VGND.n112 VGND.n84 0.146955
R663 VGND.n373 VGND.n343 0.146742
R664 VGND.n273 VGND.n272 0.146468
R665 VGND.n138 VGND.n57 0.146468
R666 VGND.n376 VGND.n340 0.146195
R667 VGND.n377 VGND.n376 0.146195
R668 VGND.n279 VGND.n278 0.146191
R669 VGND.n135 VGND.n134 0.146191
R670 VGND.n278 VGND.n277 0.145925
R671 VGND.n374 VGND.n342 0.145925
R672 VGND.n135 VGND.n60 0.145925
R673 VGND.n276 VGND.n275 0.145792
R674 VGND.n136 VGND.n59 0.145792
R675 VGND.n380 VGND.n336 0.14577
R676 VGND.n381 VGND.n335 0.14577
R677 VGND.n274 VGND.n44 0.145661
R678 VGND.n137 VGND.n58 0.145661
R679 VGND.n379 VGND.n337 0.145634
R680 VGND.n114 VGND.n82 0.145573
R681 VGND.n378 VGND.n338 0.1455
R682 VGND.n115 VGND.n81 0.145428
R683 VGND.n282 VGND.n41 0.145368
R684 VGND.n377 VGND.n339 0.145368
R685 VGND.n132 VGND.n63 0.145368
R686 VGND.n116 VGND.n80 0.145284
R687 VGND.n279 VGND.n42 0.145108
R688 VGND.n134 VGND.n61 0.145108
R689 VGND.n300 VGND.n35 0.144866
R690 VGND.n288 VGND.n39 0.144795
R691 VGND.n128 VGND.n67 0.144795
R692 VGND.n378 VGND.n377 0.144667
R693 VGND.n113 VGND.n83 0.144661
R694 VGND.n284 VGND.n283 0.14454
R695 VGND.n131 VGND.n64 0.14454
R696 VGND.n296 VGND.n295 0.144466
R697 VGND.n294 VGND.n37 0.144336
R698 VGND.n124 VGND.n71 0.144336
R699 VGND.n281 VGND.n280 0.144291
R700 VGND.n133 VGND.n62 0.144291
R701 VGND.n117 VGND.n79 0.14425
R702 VGND.n118 VGND.n78 0.144117
R703 VGND.n303 VGND.n32 0.144117
R704 VGND.n290 VGND.n289 0.144081
R705 VGND.n291 VGND.n38 0.144081
R706 VGND.n126 VGND.n69 0.144081
R707 VGND.n127 VGND.n68 0.144081
R708 VGND.n119 VGND.n77 0.143986
R709 VGND.n302 VGND.n301 0.143986
R710 VGND.n287 VGND.n286 0.143833
R711 VGND.n129 VGND.n66 0.143833
R712 VGND.n299 VGND.n298 0.143729
R713 VGND.n285 VGND.n40 0.143712
R714 VGND.n130 VGND.n65 0.143712
R715 VGND.n297 VGND.n36 0.143603
R716 VGND.n162 VGND.n158 0.143396
R717 VGND.n293 VGND.n292 0.143357
R718 VGND.n125 VGND.n70 0.143357
R719 VGND.n379 VGND.n378 0.143343
R720 VGND.n280 VGND.n41 0.142608
R721 VGND.n133 VGND.n132 0.142608
R722 VGND.n380 VGND.n379 0.142204
R723 VGND.n280 VGND.n279 0.14174
R724 VGND.n134 VGND.n133 0.14174
R725 VGND.n383 VGND.n333 0.141228
R726 VGND.n382 VGND.n381 0.140944
R727 VGND.n381 VGND.n380 0.14022
R728 VGND.n383 VGND.n382 0.139918
R729 VGND.n284 VGND.n41 0.138984
R730 VGND.n132 VGND.n131 0.138984
R731 VGND.n286 VGND.n39 0.137868
R732 VGND.n285 VGND.n284 0.137764
R733 VGND.n286 VGND.n285 0.13669
R734 VGND.n129 VGND.n128 0.135675
R735 VGND.n131 VGND.n130 0.135449
R736 VGND.n113 VGND.n112 0.134751
R737 VGND.n130 VGND.n129 0.134458
R738 VGND.n291 VGND.n290 0.134444
R739 VGND.n292 VGND.n37 0.13348
R740 VGND.n114 VGND.n113 0.133147
R741 VGND.n127 VGND.n126 0.132395
R742 VGND.n290 VGND.n39 0.132323
R743 VGND.n128 VGND.n127 0.132323
R744 VGND.n297 VGND.n296 0.131889
R745 VGND.n302 VGND.n35 0.131852
R746 VGND.n117 VGND.n116 0.13184
R747 VGND.n303 VGND.n302 0.131755
R748 VGND.n115 VGND.n114 0.131611
R749 VGND.n298 VGND.n35 0.131576
R750 VGND.n125 VGND.n124 0.131557
R751 VGND.n292 VGND.n291 0.131307
R752 VGND.n116 VGND.n115 0.131251
R753 VGND.n296 VGND.n37 0.130509
R754 VGND.n124 VGND.n123 0.130509
R755 VGND.n118 VGND.n117 0.130342
R756 VGND.n298 VGND.n297 0.130162
R757 VGND.n119 VGND.n118 0.13011
R758 VGND.n123 VGND.n122 0.130051
R759 VGND.n126 VGND.n125 0.129353
R760 VGND.n85 VGND.n84 0.124567
R761 VGND.n163 VGND.n162 0.120292
R762 VGND.n164 VGND.n163 0.120292
R763 VGND.n164 VGND.n156 0.120292
R764 VGND.n168 VGND.n156 0.120292
R765 VGND.n169 VGND.n168 0.120292
R766 VGND.n170 VGND.n169 0.120292
R767 VGND.n170 VGND.n153 0.120292
R768 VGND.n174 VGND.n153 0.120292
R769 VGND.n175 VGND.n174 0.120292
R770 VGND.n176 VGND.n175 0.120292
R771 VGND.n176 VGND.n150 0.120292
R772 VGND.n181 VGND.n150 0.120292
R773 VGND.n182 VGND.n181 0.120292
R774 VGND.n183 VGND.n182 0.120292
R775 VGND.n183 VGND.n148 0.120292
R776 VGND.n188 VGND.n148 0.120292
R777 VGND.n230 VGND.n229 0.120292
R778 VGND.n229 VGND.n193 0.120292
R779 VGND.n225 VGND.n193 0.120292
R780 VGND.n225 VGND.n224 0.120292
R781 VGND.n224 VGND.n223 0.120292
R782 VGND.n223 VGND.n195 0.120292
R783 VGND.n219 VGND.n195 0.120292
R784 VGND.n219 VGND.n218 0.120292
R785 VGND.n218 VGND.n217 0.120292
R786 VGND.n217 VGND.n198 0.120292
R787 VGND.n199 VGND.n198 0.120292
R788 VGND.n212 VGND.n199 0.120292
R789 VGND.n212 VGND.n211 0.120292
R790 VGND.n211 VGND.n202 0.120292
R791 VGND.n207 VGND.n202 0.120292
R792 VGND.n207 VGND.n206 0.120292
R793 VGND.n206 VGND.n205 0.120292
R794 VGND.n422 VGND.n421 0.120292
R795 VGND.n423 VGND.n422 0.120292
R796 VGND.n423 VGND.n23 0.120292
R797 VGND.n427 VGND.n23 0.120292
R798 VGND.n428 VGND.n427 0.120292
R799 VGND.n429 VGND.n428 0.120292
R800 VGND.n429 VGND.n20 0.120292
R801 VGND.n433 VGND.n20 0.120292
R802 VGND.n434 VGND.n433 0.120292
R803 VGND.n435 VGND.n434 0.120292
R804 VGND.n435 VGND.n18 0.120292
R805 VGND.n441 VGND.n18 0.120292
R806 VGND.n442 VGND.n441 0.120292
R807 VGND.n443 VGND.n442 0.120292
R808 VGND.n443 VGND.n16 0.120292
R809 VGND.n123 VGND.n72 0.115155
R810 VGND.n243 VGND.n55 0.110794
R811 VGND.n96 VGND.n95 0.110004
R812 VGND.n120 VGND.n76 0.109215
R813 VGND.n95 VGND.n94 0.108082
R814 VGND.n94 VGND.n93 0.105175
R815 VGND.n305 VGND.n32 0.105059
R816 VGND.n98 VGND.n96 0.104833
R817 VGND.n111 VGND.n85 0.104045
R818 VGND.n93 VGND.n92 0.1015
R819 VGND.n92 VGND.n91 0.0997064
R820 VGND VGND.n230 0.0981562
R821 VGND.n421 VGND 0.0981562
R822 VGND.n91 VGND.n90 0.097941
R823 VGND.n90 VGND.n89 0.0952266
R824 VGND.n76 VGND.n73 0.0946901
R825 VGND.n89 VGND.n88 0.0925543
R826 VGND.n460 VGND.n7 0.0910095
R827 VGND.n88 VGND.n87 0.0892405
R828 VGND.n87 VGND.n86 0.0876212
R829 VGND.n8 VGND.n7 0.0867209
R830 VGND.n457 VGND.n6 0.0867069
R831 VGND.n86 VGND.n85 0.0860263
R832 VGND.n112 VGND.n111 0.0819653
R833 VGND.n84 VGND.n83 0.0807239
R834 VGND.n122 VGND.n121 0.0803467
R835 VGND.n459 VGND.n6 0.0798478
R836 VGND.n458 VGND.n8 0.0787609
R837 VGND.n457 VGND.n456 0.0782778
R838 VGND.n97 VGND.n9 0.0776277
R839 VGND.n83 VGND.n82 0.0771423
R840 VGND.n82 VGND.n81 0.0762299
R841 VGND.n158 VGND 0.0758148
R842 VGND.n81 VGND.n80 0.0738696
R843 VGND.n97 VGND.n7 0.0721983
R844 VGND.n246 VGND.n54 0.0721201
R845 VGND.n461 VGND.n460 0.0720511
R846 VGND.n80 VGND.n79 0.0715432
R847 VGND.n79 VGND.n78 0.0701429
R848 VGND.n121 VGND.n120 0.0683371
R849 VGND.n78 VGND.n77 0.0678759
R850 VGND.n301 VGND.n32 0.0678759
R851 VGND.n72 VGND.n71 0.0675348
R852 VGND.n77 VGND.n76 0.0656408
R853 VGND.n301 VGND.n300 0.0656408
R854 VGND.n300 VGND.n299 0.0638803
R855 VGND.n299 VGND.n36 0.0621319
R856 VGND VGND.n188 0.0603958
R857 VGND.n189 VGND 0.0603958
R858 VGND.n190 VGND 0.0603958
R859 VGND.n231 VGND 0.0603958
R860 VGND.n205 VGND 0.0603958
R861 VGND.n415 VGND 0.0603958
R862 VGND.n416 VGND 0.0603958
R863 VGND.n417 VGND 0.0603958
R864 VGND.n295 VGND.n36 0.0591207
R865 VGND.n98 VGND.n97 0.0590106
R866 VGND.n295 VGND.n294 0.0582586
R867 VGND.n240 VGND 0.05675
R868 VGND.n307 VGND 0.05675
R869 VGND.n140 VGND 0.05675
R870 VGND.n34 VGND 0.05675
R871 VGND.n5 VGND 0.05675
R872 VGND.n4 VGND 0.05675
R873 VGND.n401 VGND 0.05675
R874 VGND.n3 VGND 0.05675
R875 VGND.n455 VGND 0.05675
R876 VGND.n75 VGND 0.05675
R877 VGND.n144 VGND 0.05675
R878 VGND VGND.n468 0.05675
R879 VGND.n122 VGND.n73 0.0567284
R880 VGND.n294 VGND.n293 0.0561507
R881 VGND.n71 VGND.n70 0.0561507
R882 VGND.n293 VGND.n38 0.0549218
R883 VGND.n70 VGND.n69 0.0549218
R884 VGND.n334 VGND.n333 0.0533169
R885 VGND.n289 VGND.n38 0.0520203
R886 VGND.n69 VGND.n68 0.0520203
R887 VGND.n289 VGND.n288 0.0511757
R888 VGND.n68 VGND.n67 0.0511757
R889 VGND.n387 VGND.n333 0.0509967
R890 VGND.n335 VGND.n334 0.0486419
R891 VGND.n288 VGND.n287 0.0483188
R892 VGND.n67 VGND.n66 0.0483188
R893 VGND.n336 VGND.n335 0.0477973
R894 VGND.n287 VGND.n40 0.0471667
R895 VGND.n66 VGND.n65 0.0471667
R896 VGND.n337 VGND.n336 0.045802
R897 VGND.n283 VGND.n40 0.045202
R898 VGND.n65 VGND.n64 0.045202
R899 VGND.n338 VGND.n337 0.0438333
R900 VGND.n283 VGND.n282 0.0435464
R901 VGND.n64 VGND.n63 0.0435464
R902 VGND.n282 VGND.n281 0.0418907
R903 VGND.n339 VGND.n338 0.0418907
R904 VGND.n63 VGND.n62 0.0418907
R905 VGND.n340 VGND.n339 0.0410629
R906 VGND.n458 VGND.n457 0.0407778
R907 VGND.n245 VGND.n244 0.0407077
R908 VGND.n281 VGND.n42 0.0405327
R909 VGND.n62 VGND.n61 0.0405327
R910 VGND.n341 VGND.n340 0.0385795
R911 VGND.n277 VGND.n42 0.0380817
R912 VGND.n61 VGND.n60 0.0380817
R913 VGND.n277 VGND.n276 0.0364477
R914 VGND.n342 VGND.n341 0.0364477
R915 VGND.n60 VGND.n59 0.0364477
R916 VGND.n343 VGND.n342 0.0356307
R917 VGND.n276 VGND.n44 0.0354026
R918 VGND.n59 VGND.n58 0.0354026
R919 VGND VGND.n189 0.0343542
R920 VGND VGND.n190 0.0343542
R921 VGND VGND.n415 0.0343542
R922 VGND VGND.n416 0.0343542
R923 VGND.n304 VGND.n303 0.0341879
R924 VGND.n344 VGND.n343 0.0331797
R925 VGND.n272 VGND.n44 0.0327581
R926 VGND.n58 VGND.n57 0.0327581
R927 VGND.n345 VGND.n344 0.0321558
R928 VGND.n272 VGND.n271 0.0319516
R929 VGND.n57 VGND.n56 0.0319516
R930 VGND.n73 VGND.n72 0.0307768
R931 VGND.n271 VGND.n270 0.0303387
R932 VGND.n346 VGND.n345 0.0303387
R933 VGND.n244 VGND.n56 0.0303387
R934 VGND.n456 VGND.n9 0.0297553
R935 VGND.n387 VGND.n386 0.0292963
R936 VGND.n466 VGND.n1 0.0288333
R937 VGND.n467 VGND.n466 0.0288333
R938 VGND.n347 VGND.n346 0.0279194
R939 VGND.n270 VGND.n46 0.0277436
R940 VGND.n348 VGND.n347 0.0271129
R941 VGND.n266 VGND.n46 0.0269423
R942 VGND.n349 VGND.n348 0.0253397
R943 VGND.n266 VGND.n265 0.0251815
R944 VGND.n350 VGND.n349 0.0237372
R945 VGND.n265 VGND.n264 0.0235892
R946 VGND.n231 VGND 0.0226354
R947 VGND.n417 VGND 0.0226354
R948 VGND.n264 VGND.n48 0.0219968
R949 VGND.n351 VGND.n350 0.0219968
R950 VGND.n260 VGND.n48 0.0204045
R951 VGND.n260 VGND.n259 0.0186962
R952 VGND.n275 VGND.n43 0.0175455
R953 VGND.n259 VGND.n258 0.0171139
R954 VGND.n258 VGND.n50 0.0154371
R955 VGND.n243 VGND.n242 0.0141218
R956 VGND.n254 VGND.n50 0.0139494
R957 VGND.n459 VGND.n458 0.0135435
R958 VGND.n254 VGND.n253 0.0122925
R959 VGND.n253 VGND.n252 0.00993396
R960 VGND.n365 VGND.n351 0.00918938
R961 VGND.n252 VGND.n52 0.0091478
R962 VGND.n54 VGND.n52 0.00757547
R963 VGND.n249 VGND.n248 0.00689301
R964 VGND.n465 VGND.n464 0.0011075
R965 VDPWR.n1 VDPWR.t13 738.801
R966 VDPWR.n1 VDPWR.t12 707.519
R967 VDPWR.n84 VDPWR.t63 667.734
R968 VDPWR.n52 VDPWR.t41 667.734
R969 VDPWR.n124 VDPWR.t31 667.734
R970 VDPWR.n99 VDPWR.t51 666.677
R971 VDPWR.n38 VDPWR.t59 666.677
R972 VDPWR.n4 VDPWR.t19 666.677
R973 VDPWR.t60 VDPWR.t30 624.456
R974 VDPWR.t40 VDPWR.t22 624.456
R975 VDPWR.t62 VDPWR.t24 624.456
R976 VDPWR.n102 VDPWR.n101 604.394
R977 VDPWR.n33 VDPWR.n32 604.394
R978 VDPWR.n142 VDPWR.n141 604.394
R979 VDPWR.t18 VDPWR.t52 556.386
R980 VDPWR.t32 VDPWR.t34 556.386
R981 VDPWR.t44 VDPWR.t58 556.386
R982 VDPWR.t36 VDPWR.t38 556.386
R983 VDPWR.t47 VDPWR.t50 556.386
R984 VDPWR.t66 VDPWR.t64 556.386
R985 VDPWR.n17 VDPWR.t68 414.33
R986 VDPWR.t0 VDPWR.n108 414.33
R987 VDPWR.t2 VDPWR.t6 390.654
R988 VDPWR.t72 VDPWR.t26 390.654
R989 VDPWR.t16 VDPWR.t28 390.654
R990 VDPWR.t30 VDPWR.t9 337.384
R991 VDPWR.t70 VDPWR.t40 337.384
R992 VDPWR.t56 VDPWR.t62 337.384
R993 VDPWR.n82 VDPWR.n72 333.348
R994 VDPWR.n54 VDPWR.n24 333.348
R995 VDPWR.n122 VDPWR.n12 333.348
R996 VDPWR.n68 VDPWR.n67 320.976
R997 VDPWR.n45 VDPWR.n28 320.976
R998 VDPWR.n9 VDPWR.n8 320.976
R999 VDPWR.t6 VDPWR.t55 304.829
R1000 VDPWR.t42 VDPWR.t72 304.829
R1001 VDPWR.t49 VDPWR.t16 304.829
R1002 VDPWR.t68 VDPWR.t32 287.072
R1003 VDPWR.t38 VDPWR.t0 287.072
R1004 VDPWR.t64 VDPWR.t4 287.072
R1005 VDPWR.t55 VDPWR.t8 281.154
R1006 VDPWR.t54 VDPWR.t2 281.154
R1007 VDPWR.t71 VDPWR.t42 281.154
R1008 VDPWR.t26 VDPWR.t43 281.154
R1009 VDPWR.t57 VDPWR.t49 281.154
R1010 VDPWR.t28 VDPWR.t46 281.154
R1011 VDPWR.n109 VDPWR.n17 272.274
R1012 VDPWR.n109 VDPWR 272.274
R1013 VDPWR.n108 VDPWR.n107 272.274
R1014 VDPWR.n107 VDPWR 272.274
R1015 VDPWR.t8 VDPWR.t18 251.559
R1016 VDPWR.t58 VDPWR.t71 251.559
R1017 VDPWR.t50 VDPWR.t57 251.559
R1018 VDPWR.t52 VDPWR.t20 248.599
R1019 VDPWR.t9 VDPWR.t54 248.599
R1020 VDPWR.t34 VDPWR.t60 248.599
R1021 VDPWR.t14 VDPWR.t44 248.599
R1022 VDPWR.t43 VDPWR.t70 248.599
R1023 VDPWR.t22 VDPWR.t36 248.599
R1024 VDPWR.t10 VDPWR.t47 248.599
R1025 VDPWR.t46 VDPWR.t56 248.599
R1026 VDPWR.t24 VDPWR.t66 248.599
R1027 VDPWR.n76 VDPWR.n75 240.522
R1028 VDPWR.n60 VDPWR.n21 240.522
R1029 VDPWR.n116 VDPWR.n115 240.522
R1030 VDPWR.n107 VDPWR.n106 213.119
R1031 VDPWR.n108 VDPWR.n18 213.119
R1032 VDPWR.n110 VDPWR.n109 213.119
R1033 VDPWR.n17 VDPWR.n15 213.119
R1034 VDPWR.n67 VDPWR.t17 113.98
R1035 VDPWR.n28 VDPWR.t73 113.98
R1036 VDPWR.n8 VDPWR.t7 113.98
R1037 VDPWR.t20 VDPWR 91.745
R1038 VDPWR VDPWR.t14 91.745
R1039 VDPWR VDPWR.t10 91.745
R1040 VDPWR.n75 VDPWR.t65 61.9872
R1041 VDPWR.n21 VDPWR.t39 61.9872
R1042 VDPWR.n115 VDPWR.t33 61.9872
R1043 VDPWR.n101 VDPWR.t11 41.5552
R1044 VDPWR.n101 VDPWR.t48 41.5552
R1045 VDPWR.n32 VDPWR.t15 41.5552
R1046 VDPWR.n32 VDPWR.t45 41.5552
R1047 VDPWR.n141 VDPWR.t21 41.5552
R1048 VDPWR.n141 VDPWR.t53 41.5552
R1049 VDPWR.n67 VDPWR.t29 35.4605
R1050 VDPWR.n28 VDPWR.t27 35.4605
R1051 VDPWR.n8 VDPWR.t3 35.4605
R1052 VDPWR.n81 VDPWR.n73 34.6358
R1053 VDPWR.n77 VDPWR.n73 34.6358
R1054 VDPWR.n95 VDPWR.n65 34.6358
R1055 VDPWR.n95 VDPWR.n94 34.6358
R1056 VDPWR.n94 VDPWR.n93 34.6358
R1057 VDPWR.n90 VDPWR.n89 34.6358
R1058 VDPWR.n89 VDPWR.n88 34.6358
R1059 VDPWR.n88 VDPWR.n70 34.6358
R1060 VDPWR.n55 VDPWR.n22 34.6358
R1061 VDPWR.n59 VDPWR.n22 34.6358
R1062 VDPWR.n40 VDPWR.n39 34.6358
R1063 VDPWR.n40 VDPWR.n29 34.6358
R1064 VDPWR.n44 VDPWR.n29 34.6358
R1065 VDPWR.n47 VDPWR.n46 34.6358
R1066 VDPWR.n47 VDPWR.n26 34.6358
R1067 VDPWR.n51 VDPWR.n26 34.6358
R1068 VDPWR.n121 VDPWR.n13 34.6358
R1069 VDPWR.n117 VDPWR.n13 34.6358
R1070 VDPWR.n136 VDPWR.n135 34.6358
R1071 VDPWR.n135 VDPWR.n134 34.6358
R1072 VDPWR.n134 VDPWR.n6 34.6358
R1073 VDPWR.n130 VDPWR.n129 34.6358
R1074 VDPWR.n129 VDPWR.n128 34.6358
R1075 VDPWR.n128 VDPWR.n10 34.6358
R1076 VDPWR.n83 VDPWR.n82 32.0005
R1077 VDPWR.n54 VDPWR.n53 32.0005
R1078 VDPWR.n123 VDPWR.n122 32.0005
R1079 VDPWR.n143 VDPWR.n142 30.7593
R1080 VDPWR.n84 VDPWR.n83 30.4946
R1081 VDPWR.n53 VDPWR.n52 30.4946
R1082 VDPWR.n124 VDPWR.n123 30.4946
R1083 VDPWR.n75 VDPWR.t5 30.1692
R1084 VDPWR.n21 VDPWR.t1 30.1692
R1085 VDPWR.n115 VDPWR.t69 30.1692
R1086 VDPWR.n99 VDPWR.n65 27.4829
R1087 VDPWR.n61 VDPWR.n60 27.4829
R1088 VDPWR.n39 VDPWR.n38 27.4829
R1089 VDPWR.n116 VDPWR.n114 27.4829
R1090 VDPWR.n136 VDPWR.n4 27.4829
R1091 VDPWR.n72 VDPWR.t25 26.5955
R1092 VDPWR.n72 VDPWR.t67 26.5955
R1093 VDPWR.n24 VDPWR.t23 26.5955
R1094 VDPWR.n24 VDPWR.t37 26.5955
R1095 VDPWR.n12 VDPWR.t61 26.5955
R1096 VDPWR.n12 VDPWR.t35 26.5955
R1097 VDPWR.n77 VDPWR.n76 25.6005
R1098 VDPWR.n60 VDPWR.n59 25.6005
R1099 VDPWR.n117 VDPWR.n116 25.6005
R1100 VDPWR.n106 VDPWR.n19 23.7181
R1101 VDPWR.n61 VDPWR.n18 23.7181
R1102 VDPWR.n110 VDPWR.n16 23.7181
R1103 VDPWR.n114 VDPWR.n15 23.7181
R1104 VDPWR.n102 VDPWR.n100 22.9652
R1105 VDPWR.n37 VDPWR.n33 22.9652
R1106 VDPWR.n142 VDPWR.n140 22.9652
R1107 VDPWR.n100 VDPWR.n99 21.8358
R1108 VDPWR.n38 VDPWR.n37 21.8358
R1109 VDPWR.n140 VDPWR.n4 21.8358
R1110 VDPWR.n102 VDPWR.n19 21.4593
R1111 VDPWR.n33 VDPWR.n16 21.4593
R1112 VDPWR.n93 VDPWR.n68 18.4476
R1113 VDPWR.n45 VDPWR.n44 18.4476
R1114 VDPWR.n9 VDPWR.n6 18.4476
R1115 VDPWR.n90 VDPWR.n68 16.1887
R1116 VDPWR.n46 VDPWR.n45 16.1887
R1117 VDPWR.n130 VDPWR.n9 16.1887
R1118 VDPWR.n84 VDPWR.n70 15.0593
R1119 VDPWR.n52 VDPWR.n51 15.0593
R1120 VDPWR.n124 VDPWR.n10 15.0593
R1121 VDPWR.n2 VDPWR.n1 13.3223
R1122 VDPWR.n106 VDPWR.n18 12.8005
R1123 VDPWR.n110 VDPWR.n15 12.8005
R1124 VDPWR.n3 VDPWR 9.73982
R1125 VDPWR.n143 VDPWR.n3 9.61724
R1126 VDPWR.n142 VDPWR.n0 9.3005
R1127 VDPWR.n140 VDPWR.n139 9.3005
R1128 VDPWR.n138 VDPWR.n4 9.3005
R1129 VDPWR.n137 VDPWR.n136 9.3005
R1130 VDPWR.n135 VDPWR.n5 9.3005
R1131 VDPWR.n134 VDPWR.n133 9.3005
R1132 VDPWR.n132 VDPWR.n6 9.3005
R1133 VDPWR.n131 VDPWR.n130 9.3005
R1134 VDPWR.n129 VDPWR.n7 9.3005
R1135 VDPWR.n128 VDPWR.n127 9.3005
R1136 VDPWR.n126 VDPWR.n10 9.3005
R1137 VDPWR.n125 VDPWR.n124 9.3005
R1138 VDPWR.n123 VDPWR.n11 9.3005
R1139 VDPWR.n121 VDPWR.n120 9.3005
R1140 VDPWR.n119 VDPWR.n13 9.3005
R1141 VDPWR.n118 VDPWR.n117 9.3005
R1142 VDPWR.n116 VDPWR.n14 9.3005
R1143 VDPWR.n114 VDPWR.n113 9.3005
R1144 VDPWR.n112 VDPWR.n15 9.3005
R1145 VDPWR.n111 VDPWR.n110 9.3005
R1146 VDPWR.n34 VDPWR.n16 9.3005
R1147 VDPWR.n35 VDPWR.n33 9.3005
R1148 VDPWR.n37 VDPWR.n36 9.3005
R1149 VDPWR.n38 VDPWR.n31 9.3005
R1150 VDPWR.n39 VDPWR.n30 9.3005
R1151 VDPWR.n41 VDPWR.n40 9.3005
R1152 VDPWR.n42 VDPWR.n29 9.3005
R1153 VDPWR.n44 VDPWR.n43 9.3005
R1154 VDPWR.n46 VDPWR.n27 9.3005
R1155 VDPWR.n48 VDPWR.n47 9.3005
R1156 VDPWR.n49 VDPWR.n26 9.3005
R1157 VDPWR.n51 VDPWR.n50 9.3005
R1158 VDPWR.n52 VDPWR.n25 9.3005
R1159 VDPWR.n53 VDPWR.n23 9.3005
R1160 VDPWR.n56 VDPWR.n55 9.3005
R1161 VDPWR.n57 VDPWR.n22 9.3005
R1162 VDPWR.n59 VDPWR.n58 9.3005
R1163 VDPWR.n60 VDPWR.n20 9.3005
R1164 VDPWR.n62 VDPWR.n61 9.3005
R1165 VDPWR.n63 VDPWR.n18 9.3005
R1166 VDPWR.n106 VDPWR.n105 9.3005
R1167 VDPWR.n104 VDPWR.n19 9.3005
R1168 VDPWR.n103 VDPWR.n102 9.3005
R1169 VDPWR.n100 VDPWR.n64 9.3005
R1170 VDPWR.n99 VDPWR.n98 9.3005
R1171 VDPWR.n97 VDPWR.n65 9.3005
R1172 VDPWR.n96 VDPWR.n95 9.3005
R1173 VDPWR.n94 VDPWR.n66 9.3005
R1174 VDPWR.n93 VDPWR.n92 9.3005
R1175 VDPWR.n91 VDPWR.n90 9.3005
R1176 VDPWR.n89 VDPWR.n69 9.3005
R1177 VDPWR.n88 VDPWR.n87 9.3005
R1178 VDPWR.n86 VDPWR.n70 9.3005
R1179 VDPWR.n85 VDPWR.n84 9.3005
R1180 VDPWR.n83 VDPWR.n71 9.3005
R1181 VDPWR.n81 VDPWR.n80 9.3005
R1182 VDPWR.n79 VDPWR.n73 9.3005
R1183 VDPWR.n78 VDPWR.n77 9.3005
R1184 VDPWR.n3 VDPWR.n2 8.39487
R1185 VDPWR.n76 VDPWR.n74 7.4049
R1186 VDPWR.n82 VDPWR.n81 2.63579
R1187 VDPWR.n55 VDPWR.n54 2.63579
R1188 VDPWR.n122 VDPWR.n121 2.63579
R1189 VDPWR.n74 VDPWR 0.156264
R1190 VDPWR.n78 VDPWR.n74 0.144904
R1191 VDPWR.n139 VDPWR.n0 0.120292
R1192 VDPWR.n139 VDPWR.n138 0.120292
R1193 VDPWR.n138 VDPWR.n137 0.120292
R1194 VDPWR.n137 VDPWR.n5 0.120292
R1195 VDPWR.n133 VDPWR.n5 0.120292
R1196 VDPWR.n133 VDPWR.n132 0.120292
R1197 VDPWR.n132 VDPWR.n131 0.120292
R1198 VDPWR.n131 VDPWR.n7 0.120292
R1199 VDPWR.n127 VDPWR.n7 0.120292
R1200 VDPWR.n127 VDPWR.n126 0.120292
R1201 VDPWR.n126 VDPWR.n125 0.120292
R1202 VDPWR.n125 VDPWR.n11 0.120292
R1203 VDPWR.n120 VDPWR.n11 0.120292
R1204 VDPWR.n120 VDPWR.n119 0.120292
R1205 VDPWR.n119 VDPWR.n118 0.120292
R1206 VDPWR.n118 VDPWR.n14 0.120292
R1207 VDPWR.n113 VDPWR.n14 0.120292
R1208 VDPWR.n36 VDPWR.n35 0.120292
R1209 VDPWR.n36 VDPWR.n31 0.120292
R1210 VDPWR.n31 VDPWR.n30 0.120292
R1211 VDPWR.n41 VDPWR.n30 0.120292
R1212 VDPWR.n42 VDPWR.n41 0.120292
R1213 VDPWR.n43 VDPWR.n42 0.120292
R1214 VDPWR.n43 VDPWR.n27 0.120292
R1215 VDPWR.n48 VDPWR.n27 0.120292
R1216 VDPWR.n49 VDPWR.n48 0.120292
R1217 VDPWR.n50 VDPWR.n49 0.120292
R1218 VDPWR.n50 VDPWR.n25 0.120292
R1219 VDPWR.n25 VDPWR.n23 0.120292
R1220 VDPWR.n56 VDPWR.n23 0.120292
R1221 VDPWR.n57 VDPWR.n56 0.120292
R1222 VDPWR.n58 VDPWR.n57 0.120292
R1223 VDPWR.n58 VDPWR.n20 0.120292
R1224 VDPWR.n62 VDPWR.n20 0.120292
R1225 VDPWR.n103 VDPWR.n64 0.120292
R1226 VDPWR.n98 VDPWR.n64 0.120292
R1227 VDPWR.n98 VDPWR.n97 0.120292
R1228 VDPWR.n97 VDPWR.n96 0.120292
R1229 VDPWR.n96 VDPWR.n66 0.120292
R1230 VDPWR.n92 VDPWR.n66 0.120292
R1231 VDPWR.n92 VDPWR.n91 0.120292
R1232 VDPWR.n91 VDPWR.n69 0.120292
R1233 VDPWR.n87 VDPWR.n69 0.120292
R1234 VDPWR.n87 VDPWR.n86 0.120292
R1235 VDPWR.n86 VDPWR.n85 0.120292
R1236 VDPWR.n85 VDPWR.n71 0.120292
R1237 VDPWR.n80 VDPWR.n71 0.120292
R1238 VDPWR.n80 VDPWR.n79 0.120292
R1239 VDPWR.n79 VDPWR.n78 0.120292
R1240 VDPWR VDPWR.n0 0.0981562
R1241 VDPWR.n35 VDPWR 0.0981562
R1242 VDPWR VDPWR.n103 0.0981562
R1243 VDPWR.n113 VDPWR 0.0603958
R1244 VDPWR VDPWR.n112 0.0603958
R1245 VDPWR VDPWR.n111 0.0603958
R1246 VDPWR.n34 VDPWR 0.0603958
R1247 VDPWR VDPWR.n62 0.0603958
R1248 VDPWR.n63 VDPWR 0.0603958
R1249 VDPWR.n105 VDPWR 0.0603958
R1250 VDPWR VDPWR.n104 0.0603958
R1251 VDPWR.n2 VDPWR 0.0496071
R1252 VDPWR.n112 VDPWR 0.0382604
R1253 VDPWR.n111 VDPWR 0.0382604
R1254 VDPWR VDPWR.n63 0.0382604
R1255 VDPWR.n105 VDPWR 0.0382604
R1256 VDPWR VDPWR.n34 0.0226354
R1257 VDPWR.n104 VDPWR 0.0226354
R1258 VDPWR VDPWR.n143 0.0224072
R1259 uo_out[1].n2 uo_out[1].t1 313.104
R1260 uo_out[1].n0 uo_out[1].t2 294.557
R1261 uo_out[1].t0 uo_out[1].n2 265.769
R1262 uo_out[1] uo_out[1].t0 262.318
R1263 uo_out[1].n0 uo_out[1].t3 211.01
R1264 uo_out[1].n1 uo_out[1].n0 152
R1265 uo_out[1].n5 uo_out[1] 12.6752
R1266 uo_out[1].n4 uo_out[1].n1 11.6411
R1267 uo_out[1].n4 uo_out[1].n3 9.3005
R1268 uo_out[1].n3 uo_out[1] 7.17626
R1269 uo_out[1].n3 uo_out[1].n2 4.84898
R1270 uo_out[1].n5 uo_out[1].n4 4.5029
R1271 uo_out[1].n1 uo_out[1] 1.37896
R1272 uo_out[1] uo_out[1].n5 0.0730806
R1273 uo_out[3].n0 uo_out[3].t1 313.104
R1274 uo_out[3].t0 uo_out[3].n0 265.769
R1275 uo_out[3] uo_out[3].t0 262.318
R1276 uo_out[3].n2 uo_out[3] 19.5328
R1277 uo_out[3].n2 uo_out[3].n1 13.8005
R1278 uo_out[3].n1 uo_out[3].n0 7.17626
R1279 uo_out[3].n1 uo_out[3] 4.84898
R1280 uo_out[3] uo_out[3].n2 0.0529194
R1281 uo_out[0].n0 uo_out[0].t1 983.422
R1282 uo_out[0].n7 uo_out[0].t4 543.266
R1283 uo_out[0].n8 uo_out[0].t3 526.913
R1284 uo_out[0] uo_out[0].t0 455.764
R1285 uo_out[0].n8 uo_out[0].n7 420.889
R1286 uo_out[0].n1 uo_out[0].t5 294.557
R1287 uo_out[0].n1 uo_out[0].t2 211.01
R1288 uo_out[0].n2 uo_out[0].n1 152
R1289 uo_out[0].n7 uo_out[0].n6 128.114
R1290 uo_out[0] uo_out[0].n8 125.6
R1291 uo_out[0].n6 uo_out[0].n5 60.1325
R1292 uo_out[0].n5 uo_out[0].n0 19.3454
R1293 uo_out[0].n3 uo_out[0].n2 17.6405
R1294 uo_out[0].n0 uo_out[0] 10.2862
R1295 uo_out[0] uo_out[0].n6 10.0576
R1296 uo_out[0].n4 uo_out[0].n3 6.83545
R1297 uo_out[0].n2 uo_out[0] 2.01193
R1298 uo_out[0].n4 uo_out[0] 1.31337
R1299 uo_out[0].n5 uo_out[0].n4 0.3154
R1300 uo_out[0].n3 uo_out[0] 0.0793043
R1301 uo_out[2].n2 uo_out[2].t1 313.104
R1302 uo_out[2].n0 uo_out[2].t2 294.557
R1303 uo_out[2].t0 uo_out[2].n2 265.769
R1304 uo_out[2] uo_out[2].t0 262.318
R1305 uo_out[2].n0 uo_out[2].t3 211.01
R1306 uo_out[2].n1 uo_out[2].n0 152
R1307 uo_out[2].n5 uo_out[2] 16.2155
R1308 uo_out[2].n4 uo_out[2].n1 11.6311
R1309 uo_out[2].n4 uo_out[2].n3 9.3005
R1310 uo_out[2].n3 uo_out[2] 7.17626
R1311 uo_out[2].n3 uo_out[2].n2 4.84898
R1312 uo_out[2].n5 uo_out[2].n4 4.51042
R1313 uo_out[2].n1 uo_out[2] 1.37896
R1314 uo_out[2] uo_out[2].n5 0.0730806
R1315 ua[0] ua[0].t0 973.365
R1316 ua[0].n0 ua[0].t1 466.05
R1317 ua[0] ua[0].n0 10.0576
R1318 ua[0].n0 ua[0] 7.17609
C0 m3_10182_17306# m4_10182_17306# 47.1973f
C1 m2_14954_11178# m1_14954_11178# 2.03601f
C2 m1_22770_17310# m2_22770_17310# 2.03601f
C3 m1_7076_31008# m2_7076_31008# 2.03601f
C4 m1_23290_29794# m2_23290_29794# 2.03601f
C5 m1_3616_22186# m2_3616_22186# 2.03601f
C6 m1_6556_16396# m2_6556_16396# 2.03601f
C7 m1_6556_14476# m2_6556_14476# 2.03601f
C8 VDPWR uo_out[0] 2.54419f
C9 m2_11864_11410# m1_11864_11410# 2.03601f
C10 m1_25498_23336# m2_25498_23336# 2.03601f
C11 m2_23290_27874# m1_23290_27874# 2.03601f
C12 m2_8978_14462# m1_8978_14462# 2.03601f
C13 m2_18496_31696# m1_18496_31696# 2.03601f
C14 m1_11508_25704# m2_11508_25704# 0.11049p
C15 m2_24714_24800# m1_24714_24800# 2.03601f
C16 m2_17976_11868# m1_17976_11868# 2.03601f
C17 m1_7588_42050# m2_7588_42050# 2.03601f
C18 m2_8978_12542# m1_8978_12542# 2.03601f
C19 m2_5328_28848# m1_5328_28848# 2.03601f
C20 m1_25498_21416# m2_25498_21416# 2.03601f
C21 m3_11508_25704# m2_11508_25704# 71.142296f
C22 m3_10182_17306# m2_10182_17306# 48.4105f
C23 m2_17976_13788# m1_17976_13788# 2.03601f
C24 m2_11864_13330# m1_11864_13330# 2.03601f
C25 m1_4708_16904# m2_4708_16904# 2.03601f
C26 m2_15474_34306# m1_15474_34306# 2.03601f
C27 m1_20662_15338# m2_20662_15338# 2.03601f
C28 m4_11508_25704# m3_11508_25704# 69.3594f
C29 m2_24658_17974# m1_24658_17974# 2.03601f
C30 m2_14954_13098# m1_14954_13098# 2.03601f
C31 m2_12384_32154# m1_12384_32154# 2.03601f
C32 m2_9328_42110# m1_9328_42110# 2.03601f
C33 m1_7076_29088# m2_7076_29088# 2.03601f
C34 VDPWR VAPWR 19.2978f
C35 m2_21182_32066# m1_21182_32066# 2.03601f
C36 m2_5328_26928# m1_5328_26928# 2.03601f
C37 m2_22770_15390# m1_22770_15390# 2.03601f
C38 m2_3616_20266# m1_3616_20266# 2.03601f
C39 m2_12384_34074# m1_12384_34074# 2.03601f
C40 m2_4416_25486# m1_4416_25486# 2.03601f
C41 m1_9500_32942# m2_9500_32942# 2.03601f
C42 m2_25922_1160# m1_25922_1160# 2.03601f
C43 m1_9500_31022# m2_9500_31022# 2.03601f
C44 m2_24658_19894# m1_24658_19894# 2.03601f
C45 m2_4416_23566# m1_4416_23566# 2.03601f
C46 m2_18496_33616# m1_18496_33616# 2.03601f
C47 m2_20662_13418# m1_20662_13418# 2.03601f
C48 m1_27662_1160# m2_27662_1160# 2.03601f
C49 m1_10182_17306# m2_10182_17306# 75.185295f
C50 m2_24714_26720# m1_24714_26720# 2.03601f
C51 m1_4708_18824# m2_4708_18824# 2.03601f
C52 m2_21182_30146# m1_21182_30146# 2.03601f
C53 m2_15474_32386# m1_15474_32386# 2.03601f
C54 ua[0] VGND 1.7181f
C55 uo_out[0] VGND 29.287344f
C56 uo_out[3] VGND 1.78221f
C57 VAPWR VGND 0.158964p
C58 VDPWR VGND 52.20074f
C59 m4_10182_17306# VGND 9.38538f $ **FLOATING
C60 m4_11508_25704# VGND 7.22411f $ **FLOATING
C61 m3_10182_17306# VGND 10.656599f $ **FLOATING
C62 m3_11508_25704# VGND 8.43615f $ **FLOATING
C63 m2_10182_17306# VGND 9.82879f $ **FLOATING
C64 m2_11508_25704# VGND 7.81967f $ **FLOATING
C65 m1_10182_17306# VGND 25.3587f $ **FLOATING
C66 m1_11508_25704# VGND 30.364098f $ **FLOATING
C67 ring_0/skullfet_inverter_16.A VGND 4.7412f
C68 ring_0/skullfet_inverter_17.A VGND 4.82913f
C69 ring_0/skullfet_inverter_15.A VGND 4.9312f
C70 ring_0/skullfet_inverter_18.A VGND 4.98339f
C71 ring_0/skullfet_inverter_14.A VGND 5.03686f
C72 ring_0/skullfet_inverter_19.A VGND 4.79856f
C73 ring_0/skullfet_inverter_13.A VGND 4.80717f
C74 ring_0/skullfet_inverter_20.A VGND 4.93069f
C75 ring_0/skullfet_inverter_12.A VGND 6.09378f
C76 ring_0/skullfet_inverter_20.Y VGND 5.87716f
C77 ring_0/skullfet_inverter_11.A VGND 5.42552f
C78 ring_0/skullfet_inverter_1.A VGND 5.68048f
C79 ring_0/skullfet_inverter_10.A VGND 5.3549f
C80 ring_0/skullfet_inverter_2.A VGND 5.93378f
C81 ring_0/skullfet_inverter_9.A VGND 4.59492f
C82 ring_0/skullfet_inverter_3.A VGND 5.00062f
C83 ring_0/skullfet_inverter_4.A VGND 5.01468f
C84 ring_0/skullfet_inverter_7.A VGND 4.92037f
C85 ring_0/skullfet_inverter_6.A VGND 4.74003f
C86 ring_0/skullfet_inverter_5.A VGND 4.83065f
C87 skullfet_level_shifter.A VGND 12.6722f
C88 VDPWR.n3 VGND 7.68187f
C89 VAPWR.n66 VGND 2.38783f
C90 VAPWR.n67 VGND 13.7198f
C91 VAPWR.n70 VGND 2.05887f
.ends

