MACRO tt_um_oscillating_bones
  CLASS BLOCK ;
  FOREIGN tt_um_oscillating_bones ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 143.830 224.760 144.130 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 146.590 224.760 146.890 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 141.070 224.760 141.370 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 138.310 224.760 138.610 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 135.550 224.760 135.850 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 132.790 224.760 133.090 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.030 224.760 130.330 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 127.270 224.760 127.570 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 124.510 224.760 124.810 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 121.750 224.760 122.050 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 118.990 224.760 119.290 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.230 224.760 116.530 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 113.470 224.760 113.770 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 110.710 224.760 111.010 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 107.950 224.760 108.250 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 105.190 224.760 105.490 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 102.430 224.760 102.730 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 99.670 224.760 99.970 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 96.910 224.760 97.210 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 49.990 224.760 50.290 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 47.230 224.760 47.530 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 44.470 224.760 44.770 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 41.710 224.760 42.010 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 38.950 224.760 39.250 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 36.190 224.760 36.490 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 33.430 224.760 33.730 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 30.670 224.760 30.970 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 72.070 224.760 72.370 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 69.310 224.760 69.610 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 66.550 224.760 66.850 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 63.790 224.760 64.090 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 61.030 224.760 61.330 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 58.270 224.760 58.570 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 55.510 224.760 55.810 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 52.750 224.760 53.050 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.399000 ;
    ANTENNADIFFAREA 12.700800 ;
    PORT
      LAYER met4 ;
        RECT 94.150 224.760 94.450 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 91.390 224.760 91.690 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 88.630 224.760 88.930 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 85.870 224.760 86.170 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 83.110 224.760 83.410 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 80.350 224.760 80.650 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 77.590 224.760 77.890 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 101.229294 ;
    PORT
      LAYER met4 ;
        RECT 74.830 224.760 75.130 225.760 ;
    END
  END uo_out[7]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 5.500 220.760 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 62.600 219.685 91.040 221.290 ;
      LAYER pwell ;
        RECT 62.795 219.165 65.560 219.395 ;
        RECT 67.100 219.165 68.010 219.385 ;
        RECT 62.795 218.485 71.525 219.165 ;
        RECT 71.545 218.570 71.975 219.355 ;
        RECT 72.005 218.570 72.435 219.355 ;
        RECT 72.455 219.165 75.220 219.395 ;
        RECT 76.760 219.165 77.670 219.385 ;
        RECT 72.455 218.485 81.185 219.165 ;
        RECT 81.205 218.570 81.635 219.355 ;
        RECT 81.665 218.570 82.095 219.355 ;
        RECT 82.115 219.165 84.880 219.395 ;
        RECT 86.420 219.165 87.330 219.385 ;
        RECT 82.115 218.485 90.845 219.165 ;
        RECT 71.215 218.295 71.385 218.485 ;
        RECT 80.875 218.295 81.045 218.485 ;
        RECT 90.535 218.295 90.705 218.485 ;
        RECT 65.140 174.850 70.340 180.000 ;
        RECT 82.970 176.190 88.170 181.340 ;
        RECT 48.500 168.320 53.700 173.470 ;
      LAYER nwell ;
        RECT 65.140 166.700 70.340 172.400 ;
        RECT 82.970 168.040 88.170 173.740 ;
      LAYER pwell ;
        RECT 100.410 172.210 105.610 177.360 ;
        RECT 34.510 157.170 39.710 162.320 ;
      LAYER nwell ;
        RECT 48.500 160.170 53.700 165.870 ;
        RECT 100.410 164.060 105.610 169.760 ;
      LAYER pwell ;
        RECT 115.890 163.260 121.090 168.410 ;
      LAYER nwell ;
        RECT 115.890 155.110 121.090 160.810 ;
        RECT 34.510 149.020 39.710 154.720 ;
      LAYER pwell ;
        RECT 128.060 150.150 133.260 155.300 ;
        RECT 24.440 142.390 29.640 147.540 ;
      LAYER nwell ;
        RECT 128.060 142.000 133.260 147.700 ;
        RECT 24.440 134.240 29.640 139.940 ;
      LAYER pwell ;
        RECT 136.070 134.040 141.270 139.190 ;
        RECT 19.420 125.300 24.620 130.450 ;
      LAYER nwell ;
        RECT 136.070 125.890 141.270 131.590 ;
        RECT 19.420 117.150 24.620 122.850 ;
      LAYER pwell ;
        RECT 138.490 116.360 143.690 121.510 ;
        RECT 19.170 107.420 24.370 112.570 ;
      LAYER nwell ;
        RECT 138.490 108.210 143.690 113.910 ;
        RECT 19.170 99.270 24.370 104.970 ;
      LAYER pwell ;
        RECT 136.070 98.680 141.270 103.830 ;
        RECT 24.690 90.330 29.890 95.480 ;
      LAYER nwell ;
        RECT 136.070 90.530 141.270 96.230 ;
        RECT 24.690 82.180 29.890 87.880 ;
      LAYER pwell ;
        RECT 128.310 82.570 133.510 87.720 ;
      LAYER nwell ;
        RECT 34.760 75.000 39.960 80.700 ;
      LAYER pwell ;
        RECT 34.760 67.400 39.960 72.550 ;
      LAYER nwell ;
        RECT 48.740 63.850 53.940 69.550 ;
        RECT 116.140 68.910 121.340 74.610 ;
        RECT 128.310 74.420 133.510 80.120 ;
      LAYER pwell ;
        RECT 48.740 56.250 53.940 61.400 ;
      LAYER nwell ;
        RECT 65.390 57.320 70.590 63.020 ;
        RECT 83.220 55.980 88.420 61.680 ;
        RECT 100.660 59.960 105.860 65.660 ;
      LAYER pwell ;
        RECT 116.140 61.310 121.340 66.460 ;
        RECT 65.390 49.720 70.590 54.870 ;
        RECT 83.220 48.380 88.420 53.530 ;
        RECT 100.660 52.360 105.860 57.510 ;
      LAYER li1 ;
        RECT 62.790 221.015 90.850 221.185 ;
        RECT 62.880 219.860 63.215 220.845 ;
        RECT 63.385 219.875 63.600 221.015 ;
        RECT 63.790 220.095 64.120 220.825 ;
        RECT 62.880 219.290 63.115 219.860 ;
        RECT 63.790 219.705 64.060 220.095 ;
        RECT 64.310 219.955 64.640 220.800 ;
        RECT 64.810 220.005 64.980 221.015 ;
        RECT 65.150 220.285 65.490 220.845 ;
        RECT 65.725 220.515 66.040 221.015 ;
        RECT 66.220 220.545 67.105 220.715 ;
        RECT 63.285 219.375 64.060 219.705 ;
        RECT 62.880 218.635 63.135 219.290 ;
        RECT 63.860 218.995 64.060 219.375 ;
        RECT 64.230 219.875 64.640 219.955 ;
        RECT 65.150 219.910 66.050 220.285 ;
        RECT 64.230 219.825 64.465 219.875 ;
        RECT 64.230 219.245 64.420 219.825 ;
        RECT 65.150 219.705 65.340 219.910 ;
        RECT 66.220 219.705 66.390 220.545 ;
        RECT 67.330 220.515 67.580 220.845 ;
        RECT 64.590 219.375 65.340 219.705 ;
        RECT 65.510 219.375 66.390 219.705 ;
        RECT 64.230 219.205 64.475 219.245 ;
        RECT 65.140 219.205 65.340 219.375 ;
        RECT 64.230 219.120 64.630 219.205 ;
        RECT 63.305 218.465 63.625 218.925 ;
        RECT 63.860 218.725 64.110 218.995 ;
        RECT 64.300 218.685 64.630 219.120 ;
        RECT 64.800 218.465 64.970 219.075 ;
        RECT 65.140 218.680 65.470 219.205 ;
        RECT 65.735 218.465 65.945 218.995 ;
        RECT 66.220 218.915 66.390 219.375 ;
        RECT 66.560 219.415 66.880 220.375 ;
        RECT 67.050 219.625 67.240 220.345 ;
        RECT 67.410 219.445 67.580 220.515 ;
        RECT 67.750 220.215 67.920 221.015 ;
        RECT 68.090 220.570 69.195 220.740 ;
        RECT 68.090 219.955 68.260 220.570 ;
        RECT 69.405 220.420 69.655 220.845 ;
        RECT 69.825 220.555 70.090 221.015 ;
        RECT 68.430 220.035 68.960 220.400 ;
        RECT 69.405 220.290 69.710 220.420 ;
        RECT 67.750 219.865 68.260 219.955 ;
        RECT 67.750 219.695 68.620 219.865 ;
        RECT 67.750 219.625 67.920 219.695 ;
        RECT 68.040 219.445 68.240 219.475 ;
        RECT 66.560 219.085 67.025 219.415 ;
        RECT 67.410 219.145 68.240 219.445 ;
        RECT 67.410 218.915 67.580 219.145 ;
        RECT 66.220 218.745 67.005 218.915 ;
        RECT 67.175 218.745 67.580 218.915 ;
        RECT 67.760 218.465 68.130 218.965 ;
        RECT 68.450 218.915 68.620 219.695 ;
        RECT 68.790 219.335 68.960 220.035 ;
        RECT 69.130 219.505 69.370 220.100 ;
        RECT 68.790 219.115 69.315 219.335 ;
        RECT 69.540 219.185 69.710 220.290 ;
        RECT 69.485 219.055 69.710 219.185 ;
        RECT 69.880 219.095 70.160 220.045 ;
        RECT 69.485 218.915 69.655 219.055 ;
        RECT 68.450 218.745 69.125 218.915 ;
        RECT 69.320 218.745 69.655 218.915 ;
        RECT 69.825 218.465 70.075 218.925 ;
        RECT 70.330 218.725 70.515 220.845 ;
        RECT 70.685 220.515 71.015 221.015 ;
        RECT 71.185 220.345 71.355 220.845 ;
        RECT 70.690 220.175 71.355 220.345 ;
        RECT 70.690 219.185 70.920 220.175 ;
        RECT 71.090 219.355 71.440 220.005 ;
        RECT 71.615 219.850 71.905 221.015 ;
        RECT 72.075 219.850 72.365 221.015 ;
        RECT 72.540 219.860 72.875 220.845 ;
        RECT 73.045 219.875 73.260 221.015 ;
        RECT 73.450 220.095 73.780 220.825 ;
        RECT 72.540 219.290 72.775 219.860 ;
        RECT 73.450 219.705 73.720 220.095 ;
        RECT 73.970 219.955 74.300 220.800 ;
        RECT 74.470 220.005 74.640 221.015 ;
        RECT 74.810 220.285 75.150 220.845 ;
        RECT 75.385 220.515 75.700 221.015 ;
        RECT 75.880 220.545 76.765 220.715 ;
        RECT 72.945 219.375 73.720 219.705 ;
        RECT 70.690 219.015 71.355 219.185 ;
        RECT 70.685 218.465 71.015 218.845 ;
        RECT 71.185 218.725 71.355 219.015 ;
        RECT 71.615 218.465 71.905 219.190 ;
        RECT 72.075 218.465 72.365 219.190 ;
        RECT 72.540 218.635 72.795 219.290 ;
        RECT 73.520 218.995 73.720 219.375 ;
        RECT 73.890 219.875 74.300 219.955 ;
        RECT 74.810 219.910 75.710 220.285 ;
        RECT 73.890 219.825 74.125 219.875 ;
        RECT 73.890 219.245 74.080 219.825 ;
        RECT 74.810 219.705 75.000 219.910 ;
        RECT 75.880 219.705 76.050 220.545 ;
        RECT 76.990 220.515 77.240 220.845 ;
        RECT 74.250 219.375 75.000 219.705 ;
        RECT 75.170 219.375 76.050 219.705 ;
        RECT 73.890 219.205 74.135 219.245 ;
        RECT 74.800 219.205 75.000 219.375 ;
        RECT 73.890 219.120 74.290 219.205 ;
        RECT 72.965 218.465 73.285 218.925 ;
        RECT 73.520 218.725 73.770 218.995 ;
        RECT 73.960 218.685 74.290 219.120 ;
        RECT 74.460 218.465 74.630 219.075 ;
        RECT 74.800 218.680 75.130 219.205 ;
        RECT 75.395 218.465 75.605 218.995 ;
        RECT 75.880 218.915 76.050 219.375 ;
        RECT 76.220 219.415 76.540 220.375 ;
        RECT 76.710 219.625 76.900 220.345 ;
        RECT 77.070 219.445 77.240 220.515 ;
        RECT 77.410 220.215 77.580 221.015 ;
        RECT 77.750 220.570 78.855 220.740 ;
        RECT 77.750 219.955 77.920 220.570 ;
        RECT 79.065 220.420 79.315 220.845 ;
        RECT 79.485 220.555 79.750 221.015 ;
        RECT 78.090 220.035 78.620 220.400 ;
        RECT 79.065 220.290 79.370 220.420 ;
        RECT 77.410 219.865 77.920 219.955 ;
        RECT 77.410 219.695 78.280 219.865 ;
        RECT 77.410 219.625 77.580 219.695 ;
        RECT 77.700 219.445 77.900 219.475 ;
        RECT 76.220 219.085 76.685 219.415 ;
        RECT 77.070 219.145 77.900 219.445 ;
        RECT 77.070 218.915 77.240 219.145 ;
        RECT 75.880 218.745 76.665 218.915 ;
        RECT 76.835 218.745 77.240 218.915 ;
        RECT 77.420 218.465 77.790 218.965 ;
        RECT 78.110 218.915 78.280 219.695 ;
        RECT 78.450 219.335 78.620 220.035 ;
        RECT 78.790 219.505 79.030 220.100 ;
        RECT 78.450 219.115 78.975 219.335 ;
        RECT 79.200 219.185 79.370 220.290 ;
        RECT 79.145 219.055 79.370 219.185 ;
        RECT 79.540 219.095 79.820 220.045 ;
        RECT 79.145 218.915 79.315 219.055 ;
        RECT 78.110 218.745 78.785 218.915 ;
        RECT 78.980 218.745 79.315 218.915 ;
        RECT 79.485 218.465 79.735 218.925 ;
        RECT 79.990 218.725 80.175 220.845 ;
        RECT 80.345 220.515 80.675 221.015 ;
        RECT 80.845 220.345 81.015 220.845 ;
        RECT 80.350 220.175 81.015 220.345 ;
        RECT 80.350 219.185 80.580 220.175 ;
        RECT 80.750 219.355 81.100 220.005 ;
        RECT 81.275 219.850 81.565 221.015 ;
        RECT 81.735 219.850 82.025 221.015 ;
        RECT 82.200 219.860 82.535 220.845 ;
        RECT 82.705 219.875 82.920 221.015 ;
        RECT 83.110 220.095 83.440 220.825 ;
        RECT 82.200 219.290 82.435 219.860 ;
        RECT 83.110 219.705 83.380 220.095 ;
        RECT 83.630 219.955 83.960 220.800 ;
        RECT 84.130 220.005 84.300 221.015 ;
        RECT 84.470 220.285 84.810 220.845 ;
        RECT 85.045 220.515 85.360 221.015 ;
        RECT 85.540 220.545 86.425 220.715 ;
        RECT 82.605 219.375 83.380 219.705 ;
        RECT 80.350 219.015 81.015 219.185 ;
        RECT 80.345 218.465 80.675 218.845 ;
        RECT 80.845 218.725 81.015 219.015 ;
        RECT 81.275 218.465 81.565 219.190 ;
        RECT 81.735 218.465 82.025 219.190 ;
        RECT 82.200 218.635 82.455 219.290 ;
        RECT 83.180 218.995 83.380 219.375 ;
        RECT 83.550 219.875 83.960 219.955 ;
        RECT 84.470 219.910 85.370 220.285 ;
        RECT 83.550 219.825 83.785 219.875 ;
        RECT 83.550 219.245 83.740 219.825 ;
        RECT 84.470 219.705 84.660 219.910 ;
        RECT 85.540 219.705 85.710 220.545 ;
        RECT 86.650 220.515 86.900 220.845 ;
        RECT 83.910 219.375 84.660 219.705 ;
        RECT 84.830 219.375 85.710 219.705 ;
        RECT 83.550 219.205 83.795 219.245 ;
        RECT 84.460 219.205 84.660 219.375 ;
        RECT 83.550 219.120 83.950 219.205 ;
        RECT 82.625 218.465 82.945 218.925 ;
        RECT 83.180 218.725 83.430 218.995 ;
        RECT 83.620 218.685 83.950 219.120 ;
        RECT 84.120 218.465 84.290 219.075 ;
        RECT 84.460 218.680 84.790 219.205 ;
        RECT 85.055 218.465 85.265 218.995 ;
        RECT 85.540 218.915 85.710 219.375 ;
        RECT 85.880 219.415 86.200 220.375 ;
        RECT 86.370 219.625 86.560 220.345 ;
        RECT 86.730 219.445 86.900 220.515 ;
        RECT 87.070 220.215 87.240 221.015 ;
        RECT 87.410 220.570 88.515 220.740 ;
        RECT 87.410 219.955 87.580 220.570 ;
        RECT 88.725 220.420 88.975 220.845 ;
        RECT 89.145 220.555 89.410 221.015 ;
        RECT 87.750 220.035 88.280 220.400 ;
        RECT 88.725 220.290 89.030 220.420 ;
        RECT 87.070 219.865 87.580 219.955 ;
        RECT 87.070 219.695 87.940 219.865 ;
        RECT 87.070 219.625 87.240 219.695 ;
        RECT 87.360 219.445 87.560 219.475 ;
        RECT 85.880 219.085 86.345 219.415 ;
        RECT 86.730 219.145 87.560 219.445 ;
        RECT 86.730 218.915 86.900 219.145 ;
        RECT 85.540 218.745 86.325 218.915 ;
        RECT 86.495 218.745 86.900 218.915 ;
        RECT 87.080 218.465 87.450 218.965 ;
        RECT 87.770 218.915 87.940 219.695 ;
        RECT 88.110 219.335 88.280 220.035 ;
        RECT 88.450 219.505 88.690 220.100 ;
        RECT 88.110 219.115 88.635 219.335 ;
        RECT 88.860 219.185 89.030 220.290 ;
        RECT 88.805 219.055 89.030 219.185 ;
        RECT 89.200 219.095 89.480 220.045 ;
        RECT 88.805 218.915 88.975 219.055 ;
        RECT 87.770 218.745 88.445 218.915 ;
        RECT 88.640 218.745 88.975 218.915 ;
        RECT 89.145 218.465 89.395 218.925 ;
        RECT 89.650 218.725 89.835 220.845 ;
        RECT 90.005 220.515 90.335 221.015 ;
        RECT 90.505 220.345 90.675 220.845 ;
        RECT 90.010 220.175 90.675 220.345 ;
        RECT 90.010 219.185 90.240 220.175 ;
        RECT 90.410 219.355 90.760 220.005 ;
        RECT 90.010 219.015 90.675 219.185 ;
        RECT 90.005 218.465 90.335 218.845 ;
        RECT 90.505 218.725 90.675 219.015 ;
        RECT 62.790 218.295 90.850 218.465 ;
        RECT 83.220 180.490 84.020 181.240 ;
        RECT 83.020 179.990 84.220 180.490 ;
        RECT 65.390 179.150 66.190 179.900 ;
        RECT 65.190 178.650 66.390 179.150 ;
        RECT 82.420 178.590 83.920 179.090 ;
        RECT 64.590 177.250 66.090 177.750 ;
        RECT 48.750 172.620 49.550 173.370 ;
        RECT 48.550 172.120 49.750 172.620 ;
        RECT 47.950 170.720 49.450 171.220 ;
        RECT 47.950 163.120 48.450 170.720 ;
        RECT 64.590 169.650 65.090 177.250 ;
        RECT 70.590 170.650 71.090 176.050 ;
        RECT 82.420 170.990 82.920 178.590 ;
        RECT 88.420 171.990 88.920 177.390 ;
        RECT 100.660 176.510 101.460 177.260 ;
        RECT 100.460 176.010 101.660 176.510 ;
        RECT 99.860 174.610 101.360 175.110 ;
        RECT 82.420 170.490 84.020 170.990 ;
        RECT 53.950 164.120 54.450 169.520 ;
        RECT 64.590 169.150 66.190 169.650 ;
        RECT 83.320 169.090 84.220 169.590 ;
        RECT 83.270 168.390 83.970 169.090 ;
        RECT 65.490 167.750 66.390 168.250 ;
        RECT 65.440 167.050 66.140 167.750 ;
        RECT 99.860 167.010 100.360 174.610 ;
        RECT 105.860 168.010 106.360 173.410 ;
        RECT 116.140 167.560 116.940 168.310 ;
        RECT 115.940 167.060 117.140 167.560 ;
        RECT 99.860 166.510 101.460 167.010 ;
        RECT 115.340 165.660 116.840 166.160 ;
        RECT 100.760 165.110 101.660 165.610 ;
        RECT 100.710 164.410 101.410 165.110 ;
        RECT 47.950 162.620 49.550 163.120 ;
        RECT 34.760 161.470 35.560 162.220 ;
        RECT 34.560 160.970 35.760 161.470 ;
        RECT 48.850 161.220 49.750 161.720 ;
        RECT 48.800 160.520 49.500 161.220 ;
        RECT 33.960 159.570 35.460 160.070 ;
        RECT 33.960 151.970 34.460 159.570 ;
        RECT 39.960 152.970 40.460 158.370 ;
        RECT 115.340 158.060 115.840 165.660 ;
        RECT 121.340 159.060 121.840 164.460 ;
        RECT 115.340 157.560 116.940 158.060 ;
        RECT 116.240 156.160 117.140 156.660 ;
        RECT 116.190 155.460 116.890 156.160 ;
        RECT 128.310 154.450 129.110 155.200 ;
        RECT 128.110 153.950 129.310 154.450 ;
        RECT 127.510 152.550 129.010 153.050 ;
        RECT 33.960 151.470 35.560 151.970 ;
        RECT 34.860 150.070 35.760 150.570 ;
        RECT 34.810 149.370 35.510 150.070 ;
        RECT 24.690 146.690 25.490 147.440 ;
        RECT 24.490 146.190 25.690 146.690 ;
        RECT 23.890 144.790 25.390 145.290 ;
        RECT 127.510 144.950 128.010 152.550 ;
        RECT 133.510 145.950 134.010 151.350 ;
        RECT 23.890 137.190 24.390 144.790 ;
        RECT 127.510 144.450 129.110 144.950 ;
        RECT 29.890 138.190 30.390 143.590 ;
        RECT 128.410 143.050 129.310 143.550 ;
        RECT 128.360 142.350 129.060 143.050 ;
        RECT 140.220 138.340 141.020 139.090 ;
        RECT 140.020 137.840 141.220 138.340 ;
        RECT 23.890 136.690 25.490 137.190 ;
        RECT 140.320 136.440 141.820 136.940 ;
        RECT 24.790 135.290 25.690 135.790 ;
        RECT 24.740 134.590 25.440 135.290 ;
        RECT 23.570 129.600 24.370 130.350 ;
        RECT 135.320 129.840 135.820 135.240 ;
        RECT 23.370 129.100 24.570 129.600 ;
        RECT 141.320 128.840 141.820 136.440 ;
        RECT 140.220 128.340 141.820 128.840 ;
        RECT 23.670 127.700 25.170 128.200 ;
        RECT 18.670 121.100 19.170 126.500 ;
        RECT 24.670 120.100 25.170 127.700 ;
        RECT 140.020 126.940 140.920 127.440 ;
        RECT 140.270 126.240 140.970 126.940 ;
        RECT 138.740 120.660 139.540 121.410 ;
        RECT 138.540 120.160 139.740 120.660 ;
        RECT 23.570 119.600 25.170 120.100 ;
        RECT 137.940 118.760 139.440 119.260 ;
        RECT 23.370 118.200 24.270 118.700 ;
        RECT 23.620 117.500 24.320 118.200 ;
        RECT 19.420 111.720 20.220 112.470 ;
        RECT 19.220 111.220 20.420 111.720 ;
        RECT 137.940 111.160 138.440 118.760 ;
        RECT 143.940 112.160 144.440 117.560 ;
        RECT 137.940 110.660 139.540 111.160 ;
        RECT 18.620 109.820 20.120 110.320 ;
        RECT 18.620 102.220 19.120 109.820 ;
        RECT 138.840 109.260 139.740 109.760 ;
        RECT 24.620 103.220 25.120 108.620 ;
        RECT 138.790 108.560 139.490 109.260 ;
        RECT 140.220 102.980 141.020 103.730 ;
        RECT 140.020 102.480 141.220 102.980 ;
        RECT 18.620 101.720 20.220 102.220 ;
        RECT 140.320 101.080 141.820 101.580 ;
        RECT 19.520 100.320 20.420 100.820 ;
        RECT 19.470 99.620 20.170 100.320 ;
        RECT 28.840 94.630 29.640 95.380 ;
        RECT 28.640 94.130 29.840 94.630 ;
        RECT 135.320 94.480 135.820 99.880 ;
        RECT 141.320 93.480 141.820 101.080 ;
        RECT 28.940 92.730 30.440 93.230 ;
        RECT 140.220 92.980 141.820 93.480 ;
        RECT 23.940 86.130 24.440 91.530 ;
        RECT 29.940 85.130 30.440 92.730 ;
        RECT 140.020 91.580 140.920 92.080 ;
        RECT 140.270 90.880 140.970 91.580 ;
        RECT 132.460 86.870 133.260 87.620 ;
        RECT 132.260 86.370 133.460 86.870 ;
        RECT 28.840 84.630 30.440 85.130 ;
        RECT 132.560 84.970 134.060 85.470 ;
        RECT 28.640 83.230 29.540 83.730 ;
        RECT 28.890 82.530 29.590 83.230 ;
        RECT 38.960 79.650 39.660 80.350 ;
        RECT 38.710 79.150 39.610 79.650 ;
        RECT 127.560 78.370 128.060 83.770 ;
        RECT 38.910 77.750 40.510 78.250 ;
        RECT 34.010 71.350 34.510 76.750 ;
        RECT 40.010 70.150 40.510 77.750 ;
        RECT 133.560 77.370 134.060 84.970 ;
        RECT 132.460 76.870 134.060 77.370 ;
        RECT 132.260 75.470 133.160 75.970 ;
        RECT 132.510 74.770 133.210 75.470 ;
        RECT 120.340 73.560 121.040 74.260 ;
        RECT 120.090 73.060 120.990 73.560 ;
        RECT 120.290 71.660 121.890 72.160 ;
        RECT 39.010 69.650 40.510 70.150 ;
        RECT 38.710 68.250 39.910 68.750 ;
        RECT 52.940 68.500 53.640 69.200 ;
        RECT 38.910 67.500 39.710 68.250 ;
        RECT 52.690 68.000 53.590 68.500 ;
        RECT 52.890 66.600 54.490 67.100 ;
        RECT 47.990 60.200 48.490 65.600 ;
        RECT 53.990 59.000 54.490 66.600 ;
        RECT 104.860 64.610 105.560 65.310 ;
        RECT 115.390 65.260 115.890 70.660 ;
        RECT 104.610 64.110 105.510 64.610 ;
        RECT 121.390 64.060 121.890 71.660 ;
        RECT 120.390 63.560 121.890 64.060 ;
        RECT 104.810 62.710 106.410 63.210 ;
        RECT 69.590 61.970 70.290 62.670 ;
        RECT 69.340 61.470 70.240 61.970 ;
        RECT 87.420 60.630 88.120 61.330 ;
        RECT 69.540 60.070 71.140 60.570 ;
        RECT 87.170 60.130 88.070 60.630 ;
        RECT 52.990 58.500 54.490 59.000 ;
        RECT 52.690 57.100 53.890 57.600 ;
        RECT 52.890 56.350 53.690 57.100 ;
        RECT 64.640 53.670 65.140 59.070 ;
        RECT 70.640 52.470 71.140 60.070 ;
        RECT 87.370 58.730 88.970 59.230 ;
        RECT 69.640 51.970 71.140 52.470 ;
        RECT 82.470 52.330 82.970 57.730 ;
        RECT 88.470 51.130 88.970 58.730 ;
        RECT 99.910 56.310 100.410 61.710 ;
        RECT 105.910 55.110 106.410 62.710 ;
        RECT 120.090 62.160 121.290 62.660 ;
        RECT 120.290 61.410 121.090 62.160 ;
        RECT 104.910 54.610 106.410 55.110 ;
        RECT 104.610 53.210 105.810 53.710 ;
        RECT 104.810 52.460 105.610 53.210 ;
        RECT 69.340 50.570 70.540 51.070 ;
        RECT 87.470 50.630 88.970 51.130 ;
        RECT 69.540 49.820 70.340 50.570 ;
        RECT 87.170 49.230 88.370 49.730 ;
        RECT 87.370 48.480 88.170 49.230 ;
      LAYER met1 ;
        RECT 90.535 221.340 92.300 221.345 ;
        RECT 62.790 220.865 92.300 221.340 ;
        RECT 62.790 220.860 90.850 220.865 ;
        RECT 67.000 220.320 67.290 220.365 ;
        RECT 68.570 220.320 68.860 220.365 ;
        RECT 70.670 220.320 70.960 220.365 ;
        RECT 67.000 220.180 70.960 220.320 ;
        RECT 67.000 220.135 67.290 220.180 ;
        RECT 68.570 220.135 68.860 220.180 ;
        RECT 70.670 220.135 70.960 220.180 ;
        RECT 76.660 220.320 76.950 220.365 ;
        RECT 78.230 220.320 78.520 220.365 ;
        RECT 80.330 220.320 80.620 220.365 ;
        RECT 76.660 220.180 80.620 220.320 ;
        RECT 76.660 220.135 76.950 220.180 ;
        RECT 78.230 220.135 78.520 220.180 ;
        RECT 80.330 220.135 80.620 220.180 ;
        RECT 86.320 220.320 86.610 220.365 ;
        RECT 87.890 220.320 88.180 220.365 ;
        RECT 89.990 220.320 90.280 220.365 ;
        RECT 86.320 220.180 90.280 220.320 ;
        RECT 86.320 220.135 86.610 220.180 ;
        RECT 87.890 220.135 88.180 220.180 ;
        RECT 89.990 220.135 90.280 220.180 ;
        RECT 62.880 219.870 63.170 220.100 ;
        RECT 66.565 219.980 66.855 220.025 ;
        RECT 69.085 219.980 69.375 220.025 ;
        RECT 70.275 219.980 70.565 220.025 ;
        RECT 62.990 219.640 63.130 219.870 ;
        RECT 66.565 219.840 70.565 219.980 ;
        RECT 72.535 219.870 72.825 220.100 ;
        RECT 76.225 219.980 76.515 220.025 ;
        RECT 78.745 219.980 79.035 220.025 ;
        RECT 79.935 219.980 80.225 220.025 ;
        RECT 66.565 219.795 66.855 219.840 ;
        RECT 69.085 219.795 69.375 219.840 ;
        RECT 70.275 219.795 70.565 219.840 ;
        RECT 69.850 219.640 70.140 219.680 ;
        RECT 62.990 219.500 70.140 219.640 ;
        RECT 69.850 219.450 70.140 219.500 ;
        RECT 71.140 219.425 71.430 219.655 ;
        RECT 72.645 219.640 72.785 219.870 ;
        RECT 76.225 219.840 80.225 219.980 ;
        RECT 82.200 219.870 82.490 220.100 ;
        RECT 85.885 219.980 86.175 220.025 ;
        RECT 88.405 219.980 88.695 220.025 ;
        RECT 89.595 219.980 89.885 220.025 ;
        RECT 76.225 219.795 76.515 219.840 ;
        RECT 78.745 219.795 79.035 219.840 ;
        RECT 79.935 219.795 80.225 219.840 ;
        RECT 79.505 219.640 79.795 219.680 ;
        RECT 72.645 219.500 79.795 219.640 ;
        RECT 79.505 219.450 79.795 219.500 ;
        RECT 80.800 219.425 81.090 219.655 ;
        RECT 82.310 219.640 82.450 219.870 ;
        RECT 85.885 219.840 89.885 219.980 ;
        RECT 90.440 219.840 90.720 219.900 ;
        RECT 85.885 219.795 86.175 219.840 ;
        RECT 88.405 219.795 88.695 219.840 ;
        RECT 89.595 219.795 89.885 219.840 ;
        RECT 89.170 219.640 89.460 219.680 ;
        RECT 82.310 219.500 89.460 219.640 ;
        RECT 89.170 219.450 89.460 219.500 ;
        RECT 90.380 219.455 90.740 219.840 ;
        RECT 64.260 218.770 64.690 219.090 ;
        RECT 71.200 219.075 71.370 219.425 ;
        RECT 73.975 219.075 74.265 219.105 ;
        RECT 71.200 219.020 74.265 219.075 ;
        RECT 80.860 219.075 81.030 219.425 ;
        RECT 90.440 219.395 90.720 219.455 ;
        RECT 83.580 219.075 83.990 219.120 ;
        RECT 71.200 218.905 74.350 219.020 ;
        RECT 80.860 218.905 83.990 219.075 ;
        RECT 73.940 218.760 74.350 218.905 ;
        RECT 83.580 218.860 83.990 218.905 ;
        RECT 61.430 218.140 90.850 218.620 ;
        RECT 84.650 180.740 86.810 181.010 ;
        RECT 82.420 180.490 82.820 180.590 ;
        RECT 82.420 180.040 83.420 180.490 ;
        RECT 84.380 180.470 86.810 180.740 ;
        RECT 83.840 179.930 87.350 180.470 ;
        RECT 66.820 179.400 68.980 179.670 ;
        RECT 64.590 179.150 64.990 179.250 ;
        RECT 64.590 178.700 65.590 179.150 ;
        RECT 66.550 179.130 68.980 179.400 ;
        RECT 66.010 178.590 69.520 179.130 ;
        RECT 83.570 178.850 87.620 179.930 ;
        RECT 65.740 177.510 69.790 178.590 ;
        RECT 83.570 178.580 84.380 178.850 ;
        RECT 83.570 178.310 84.110 178.580 ;
        RECT 65.740 177.240 66.550 177.510 ;
        RECT 65.740 176.970 66.280 177.240 ;
        RECT 66.010 176.700 66.280 176.970 ;
        RECT 67.360 176.700 68.170 177.510 ;
        RECT 68.980 177.240 69.790 177.510 ;
        RECT 83.840 178.040 84.110 178.310 ;
        RECT 85.190 178.040 86.000 178.850 ;
        RECT 86.810 178.580 87.620 178.850 ;
        RECT 87.080 178.310 87.620 178.580 ;
        RECT 87.080 178.040 87.350 178.310 ;
        RECT 83.840 177.770 84.380 178.040 ;
        RECT 84.920 177.770 86.270 178.040 ;
        RECT 86.810 177.770 87.350 178.040 ;
        RECT 83.840 177.500 85.460 177.770 ;
        RECT 85.730 177.500 87.080 177.770 ;
        RECT 69.250 176.970 69.790 177.240 ;
        RECT 84.380 177.230 85.190 177.500 ;
        RECT 86.000 177.230 87.080 177.500 ;
        RECT 69.250 176.700 69.520 176.970 ;
        RECT 66.010 176.430 66.550 176.700 ;
        RECT 67.090 176.430 68.440 176.700 ;
        RECT 68.980 176.430 69.520 176.700 ;
        RECT 84.650 176.690 86.540 177.230 ;
        RECT 102.090 176.760 104.250 177.030 ;
        RECT 66.010 176.160 67.630 176.430 ;
        RECT 67.900 176.160 69.250 176.430 ;
        RECT 83.030 176.420 83.840 176.690 ;
        RECT 84.650 176.420 84.920 176.690 ;
        RECT 85.190 176.420 85.460 176.690 ;
        RECT 85.730 176.420 86.000 176.690 ;
        RECT 86.270 176.420 86.540 176.690 ;
        RECT 87.350 176.420 88.160 176.690 ;
        RECT 99.860 176.510 100.260 176.610 ;
        RECT 66.550 175.890 67.360 176.160 ;
        RECT 68.170 175.890 69.250 176.160 ;
        RECT 66.820 175.350 68.710 175.890 ;
        RECT 82.760 175.880 84.110 176.420 ;
        RECT 87.080 175.880 88.430 176.420 ;
        RECT 99.860 176.060 100.860 176.510 ;
        RECT 101.820 176.490 104.250 176.760 ;
        RECT 101.280 175.950 104.790 176.490 ;
        RECT 83.030 175.610 84.650 175.880 ;
        RECT 86.540 175.610 88.160 175.880 ;
        RECT 65.200 175.080 66.010 175.350 ;
        RECT 66.820 175.080 67.090 175.350 ;
        RECT 67.360 175.080 67.630 175.350 ;
        RECT 67.900 175.080 68.170 175.350 ;
        RECT 68.440 175.080 68.710 175.350 ;
        RECT 69.520 175.080 70.330 175.350 ;
        RECT 76.705 175.340 82.335 175.345 ;
        RECT 83.840 175.340 84.920 175.610 ;
        RECT 86.270 175.340 87.350 175.610 ;
        RECT 64.930 174.540 66.280 175.080 ;
        RECT 69.250 174.540 70.600 175.080 ;
        RECT 76.705 174.795 82.920 175.340 ;
        RECT 84.380 175.070 85.460 175.340 ;
        RECT 85.730 175.070 86.810 175.340 ;
        RECT 88.420 175.165 89.420 175.340 ;
        RECT 65.200 174.270 66.820 174.540 ;
        RECT 68.710 174.270 70.330 174.540 ;
        RECT 66.010 174.000 67.090 174.270 ;
        RECT 68.440 174.000 69.520 174.270 ;
        RECT 64.140 173.945 65.090 174.000 ;
        RECT 58.375 173.395 65.090 173.945 ;
        RECT 66.550 173.730 67.630 174.000 ;
        RECT 67.900 173.730 68.980 174.000 ;
        RECT 70.590 173.865 71.590 174.000 ;
        RECT 76.705 173.865 77.255 174.795 ;
        RECT 81.970 174.440 82.920 174.795 ;
        RECT 84.920 174.530 86.270 175.070 ;
        RECT 88.420 174.615 97.185 175.165 ;
        RECT 84.380 174.260 85.460 174.530 ;
        RECT 85.730 174.260 86.810 174.530 ;
        RECT 88.420 174.440 89.420 174.615 ;
        RECT 83.030 173.990 84.920 174.260 ;
        RECT 86.270 173.990 88.430 174.260 ;
        RECT 50.180 172.870 52.340 173.140 ;
        RECT 47.950 172.620 48.350 172.720 ;
        RECT 47.950 172.170 48.950 172.620 ;
        RECT 49.910 172.600 52.340 172.870 ;
        RECT 49.370 172.060 52.880 172.600 ;
        RECT 49.100 170.980 53.150 172.060 ;
        RECT 49.100 170.710 49.910 170.980 ;
        RECT 49.100 170.440 49.640 170.710 ;
        RECT 49.370 170.170 49.640 170.440 ;
        RECT 50.720 170.170 51.530 170.980 ;
        RECT 52.340 170.710 53.150 170.980 ;
        RECT 52.610 170.440 53.150 170.710 ;
        RECT 52.610 170.170 52.880 170.440 ;
        RECT 49.370 169.900 49.910 170.170 ;
        RECT 50.450 169.900 51.800 170.170 ;
        RECT 52.340 169.900 52.880 170.170 ;
        RECT 49.370 169.630 50.990 169.900 ;
        RECT 51.260 169.630 52.610 169.900 ;
        RECT 49.910 169.360 50.720 169.630 ;
        RECT 51.530 169.360 52.610 169.630 ;
        RECT 50.180 168.820 52.070 169.360 ;
        RECT 48.560 168.550 49.370 168.820 ;
        RECT 50.180 168.550 50.450 168.820 ;
        RECT 50.720 168.550 50.990 168.820 ;
        RECT 51.260 168.550 51.530 168.820 ;
        RECT 51.800 168.550 52.070 168.820 ;
        RECT 52.880 168.550 53.690 168.820 ;
        RECT 48.290 168.010 49.640 168.550 ;
        RECT 52.610 168.010 53.960 168.550 ;
        RECT 48.560 167.740 50.180 168.010 ;
        RECT 52.070 167.740 53.690 168.010 ;
        RECT 49.370 167.470 50.450 167.740 ;
        RECT 51.800 167.470 52.880 167.740 ;
        RECT 47.500 167.240 48.450 167.470 ;
        RECT 43.210 166.740 48.450 167.240 ;
        RECT 49.910 167.200 50.990 167.470 ;
        RECT 51.260 167.200 52.340 167.470 ;
        RECT 53.950 167.365 54.950 167.470 ;
        RECT 58.375 167.365 58.925 173.395 ;
        RECT 64.140 173.100 65.090 173.395 ;
        RECT 67.090 173.190 68.440 173.730 ;
        RECT 70.590 173.315 77.255 173.865 ;
        RECT 82.760 173.720 84.380 173.990 ;
        RECT 86.810 173.720 88.430 173.990 ;
        RECT 82.760 173.450 83.840 173.720 ;
        RECT 87.350 173.450 88.430 173.720 ;
        RECT 66.550 172.920 67.630 173.190 ;
        RECT 67.900 172.920 68.980 173.190 ;
        RECT 70.590 173.100 71.590 173.315 ;
        RECT 82.760 173.180 83.570 173.450 ;
        RECT 87.620 173.180 88.430 173.450 ;
        RECT 65.200 172.650 67.090 172.920 ;
        RECT 68.440 172.650 70.600 172.920 ;
        RECT 83.030 172.910 83.300 173.180 ;
        RECT 84.650 172.910 84.920 173.180 ;
        RECT 85.190 172.910 85.460 173.180 ;
        RECT 85.730 172.910 86.000 173.180 ;
        RECT 86.270 172.910 86.540 173.180 ;
        RECT 87.890 172.910 88.160 173.180 ;
        RECT 64.930 172.380 66.550 172.650 ;
        RECT 68.980 172.380 70.600 172.650 ;
        RECT 64.930 172.110 66.010 172.380 ;
        RECT 69.520 172.110 70.600 172.380 ;
        RECT 84.650 172.370 86.540 172.910 ;
        RECT 64.930 171.840 65.740 172.110 ;
        RECT 69.790 171.840 70.600 172.110 ;
        RECT 84.380 172.100 85.190 172.370 ;
        RECT 86.000 172.100 87.080 172.370 ;
        RECT 65.200 171.570 65.470 171.840 ;
        RECT 66.820 171.570 67.090 171.840 ;
        RECT 67.360 171.570 67.630 171.840 ;
        RECT 67.900 171.570 68.170 171.840 ;
        RECT 68.440 171.570 68.710 171.840 ;
        RECT 70.060 171.570 70.330 171.840 ;
        RECT 83.840 171.830 85.460 172.100 ;
        RECT 85.730 171.830 87.080 172.100 ;
        RECT 66.820 171.030 68.710 171.570 ;
        RECT 83.840 171.560 84.380 171.830 ;
        RECT 84.920 171.560 86.270 171.830 ;
        RECT 86.810 171.560 87.350 171.830 ;
        RECT 83.840 171.290 84.110 171.560 ;
        RECT 66.550 170.760 67.360 171.030 ;
        RECT 68.170 170.760 69.250 171.030 ;
        RECT 66.010 170.490 67.630 170.760 ;
        RECT 67.900 170.490 69.250 170.760 ;
        RECT 83.570 171.020 84.110 171.290 ;
        RECT 83.570 170.750 84.380 171.020 ;
        RECT 85.190 170.750 86.000 171.560 ;
        RECT 87.080 171.290 87.350 171.560 ;
        RECT 87.080 171.020 87.620 171.290 ;
        RECT 86.810 170.750 87.620 171.020 ;
        RECT 66.010 170.220 66.550 170.490 ;
        RECT 67.090 170.220 68.440 170.490 ;
        RECT 68.980 170.220 69.520 170.490 ;
        RECT 66.010 169.950 66.280 170.220 ;
        RECT 65.740 169.680 66.280 169.950 ;
        RECT 65.740 169.410 66.550 169.680 ;
        RECT 67.360 169.410 68.170 170.220 ;
        RECT 69.250 169.950 69.520 170.220 ;
        RECT 69.250 169.680 69.790 169.950 ;
        RECT 68.980 169.410 69.790 169.680 ;
        RECT 83.570 169.670 87.620 170.750 ;
        RECT 96.635 171.165 97.185 174.615 ;
        RECT 101.010 174.870 105.060 175.950 ;
        RECT 101.010 174.600 101.820 174.870 ;
        RECT 101.010 174.330 101.550 174.600 ;
        RECT 101.280 174.060 101.550 174.330 ;
        RECT 102.630 174.060 103.440 174.870 ;
        RECT 104.250 174.600 105.060 174.870 ;
        RECT 104.520 174.330 105.060 174.600 ;
        RECT 104.520 174.060 104.790 174.330 ;
        RECT 101.280 173.790 101.820 174.060 ;
        RECT 102.360 173.790 103.710 174.060 ;
        RECT 104.250 173.790 104.790 174.060 ;
        RECT 101.280 173.520 102.900 173.790 ;
        RECT 103.170 173.520 104.520 173.790 ;
        RECT 101.820 173.250 102.630 173.520 ;
        RECT 103.440 173.250 104.520 173.520 ;
        RECT 102.090 172.710 103.980 173.250 ;
        RECT 100.470 172.440 101.280 172.710 ;
        RECT 102.090 172.440 102.360 172.710 ;
        RECT 102.630 172.440 102.900 172.710 ;
        RECT 103.170 172.440 103.440 172.710 ;
        RECT 103.710 172.440 103.980 172.710 ;
        RECT 104.790 172.440 105.600 172.710 ;
        RECT 100.200 171.900 101.550 172.440 ;
        RECT 104.520 171.900 105.870 172.440 ;
        RECT 100.470 171.630 102.090 171.900 ;
        RECT 103.980 171.630 105.600 171.900 ;
        RECT 101.280 171.360 102.360 171.630 ;
        RECT 103.710 171.360 104.790 171.630 ;
        RECT 99.410 171.165 100.360 171.360 ;
        RECT 96.635 170.615 100.360 171.165 ;
        RECT 101.820 171.090 102.900 171.360 ;
        RECT 103.170 171.090 104.250 171.360 ;
        RECT 105.860 171.185 106.860 171.360 ;
        RECT 99.410 170.460 100.360 170.615 ;
        RECT 102.360 170.550 103.710 171.090 ;
        RECT 105.860 170.635 110.815 171.185 ;
        RECT 101.820 170.280 102.900 170.550 ;
        RECT 103.170 170.280 104.250 170.550 ;
        RECT 105.860 170.460 106.860 170.635 ;
        RECT 100.470 170.010 102.360 170.280 ;
        RECT 103.710 170.010 105.870 170.280 ;
        RECT 100.200 169.740 101.820 170.010 ;
        RECT 104.250 169.740 105.870 170.010 ;
        RECT 65.740 168.330 69.790 169.410 ;
        RECT 82.420 169.090 83.670 169.490 ;
        RECT 83.840 169.130 87.350 169.670 ;
        RECT 100.200 169.470 101.280 169.740 ;
        RECT 104.790 169.470 105.870 169.740 ;
        RECT 100.200 169.200 101.010 169.470 ;
        RECT 105.060 169.200 105.870 169.470 ;
        RECT 82.420 168.940 82.920 169.090 ;
        RECT 84.380 168.860 86.810 169.130 ;
        RECT 100.470 168.930 100.740 169.200 ;
        RECT 102.090 168.930 102.360 169.200 ;
        RECT 102.630 168.930 102.900 169.200 ;
        RECT 103.170 168.930 103.440 169.200 ;
        RECT 103.710 168.930 103.980 169.200 ;
        RECT 105.330 168.930 105.600 169.200 ;
        RECT 84.650 168.590 86.810 168.860 ;
        RECT 102.090 168.390 103.980 168.930 ;
        RECT 64.590 167.750 65.840 168.150 ;
        RECT 66.010 167.790 69.520 168.330 ;
        RECT 101.820 168.120 102.630 168.390 ;
        RECT 103.440 168.120 104.520 168.390 ;
        RECT 101.280 167.850 102.900 168.120 ;
        RECT 103.170 167.850 104.520 168.120 ;
        RECT 64.590 167.600 65.090 167.750 ;
        RECT 66.550 167.520 68.980 167.790 ;
        RECT 36.190 161.720 38.350 161.990 ;
        RECT 33.960 161.470 34.360 161.570 ;
        RECT 33.960 161.020 34.960 161.470 ;
        RECT 35.920 161.450 38.350 161.720 ;
        RECT 35.380 160.910 38.890 161.450 ;
        RECT 35.110 159.830 39.160 160.910 ;
        RECT 35.110 159.560 35.920 159.830 ;
        RECT 35.110 159.290 35.650 159.560 ;
        RECT 35.380 159.020 35.650 159.290 ;
        RECT 36.730 159.020 37.540 159.830 ;
        RECT 38.350 159.560 39.160 159.830 ;
        RECT 38.620 159.290 39.160 159.560 ;
        RECT 38.620 159.020 38.890 159.290 ;
        RECT 35.380 158.750 35.920 159.020 ;
        RECT 36.460 158.750 37.810 159.020 ;
        RECT 38.350 158.750 38.890 159.020 ;
        RECT 35.380 158.480 37.000 158.750 ;
        RECT 37.270 158.480 38.620 158.750 ;
        RECT 35.920 158.210 36.730 158.480 ;
        RECT 37.540 158.210 38.620 158.480 ;
        RECT 36.190 157.670 38.080 158.210 ;
        RECT 34.570 157.400 35.380 157.670 ;
        RECT 36.190 157.400 36.460 157.670 ;
        RECT 36.730 157.400 37.000 157.670 ;
        RECT 37.270 157.400 37.540 157.670 ;
        RECT 37.810 157.400 38.080 157.670 ;
        RECT 38.890 157.400 39.700 157.670 ;
        RECT 34.300 156.860 35.650 157.400 ;
        RECT 38.620 156.860 39.970 157.400 ;
        RECT 34.570 156.590 36.190 156.860 ;
        RECT 38.080 156.590 39.700 156.860 ;
        RECT 35.380 156.320 36.460 156.590 ;
        RECT 37.810 156.320 38.890 156.590 ;
        RECT 33.510 156.100 34.460 156.320 ;
        RECT 30.880 155.600 34.460 156.100 ;
        RECT 35.920 156.050 37.000 156.320 ;
        RECT 37.270 156.050 38.350 156.320 ;
        RECT 39.960 156.130 40.960 156.320 ;
        RECT 43.210 156.130 43.710 166.740 ;
        RECT 47.500 166.570 48.450 166.740 ;
        RECT 50.450 166.660 51.800 167.200 ;
        RECT 53.950 166.815 58.925 167.365 ;
        RECT 66.820 167.250 68.980 167.520 ;
        RECT 101.280 167.580 101.820 167.850 ;
        RECT 102.360 167.580 103.710 167.850 ;
        RECT 104.250 167.580 104.790 167.850 ;
        RECT 101.280 167.310 101.550 167.580 ;
        RECT 101.010 167.040 101.550 167.310 ;
        RECT 49.910 166.390 50.990 166.660 ;
        RECT 51.260 166.390 52.340 166.660 ;
        RECT 53.950 166.570 54.950 166.815 ;
        RECT 101.010 166.770 101.820 167.040 ;
        RECT 102.630 166.770 103.440 167.580 ;
        RECT 104.520 167.310 104.790 167.580 ;
        RECT 104.520 167.040 105.060 167.310 ;
        RECT 104.250 166.770 105.060 167.040 ;
        RECT 48.560 166.120 50.450 166.390 ;
        RECT 51.800 166.120 53.960 166.390 ;
        RECT 48.290 165.850 49.910 166.120 ;
        RECT 52.340 165.850 53.960 166.120 ;
        RECT 48.290 165.580 49.370 165.850 ;
        RECT 52.880 165.580 53.960 165.850 ;
        RECT 101.010 165.690 105.060 166.770 ;
        RECT 48.290 165.310 49.100 165.580 ;
        RECT 53.150 165.310 53.960 165.580 ;
        RECT 48.560 165.040 48.830 165.310 ;
        RECT 50.180 165.040 50.450 165.310 ;
        RECT 50.720 165.040 50.990 165.310 ;
        RECT 51.260 165.040 51.530 165.310 ;
        RECT 51.800 165.040 52.070 165.310 ;
        RECT 53.420 165.040 53.690 165.310 ;
        RECT 99.860 165.110 101.110 165.510 ;
        RECT 101.280 165.150 104.790 165.690 ;
        RECT 50.180 164.500 52.070 165.040 ;
        RECT 99.860 164.960 100.360 165.110 ;
        RECT 101.820 164.880 104.250 165.150 ;
        RECT 102.090 164.610 104.250 164.880 ;
        RECT 49.910 164.230 50.720 164.500 ;
        RECT 51.530 164.230 52.610 164.500 ;
        RECT 49.370 163.960 50.990 164.230 ;
        RECT 51.260 163.960 52.610 164.230 ;
        RECT 49.370 163.690 49.910 163.960 ;
        RECT 50.450 163.690 51.800 163.960 ;
        RECT 52.340 163.690 52.880 163.960 ;
        RECT 49.370 163.420 49.640 163.690 ;
        RECT 49.100 163.150 49.640 163.420 ;
        RECT 49.100 162.880 49.910 163.150 ;
        RECT 50.720 162.880 51.530 163.690 ;
        RECT 52.610 163.420 52.880 163.690 ;
        RECT 52.610 163.150 53.150 163.420 ;
        RECT 52.340 162.880 53.150 163.150 ;
        RECT 49.100 161.800 53.150 162.880 ;
        RECT 110.265 162.135 110.815 170.635 ;
        RECT 117.570 167.810 119.730 168.080 ;
        RECT 115.340 167.560 115.740 167.660 ;
        RECT 115.340 167.110 116.340 167.560 ;
        RECT 117.300 167.540 119.730 167.810 ;
        RECT 116.760 167.000 120.270 167.540 ;
        RECT 116.490 165.920 120.540 167.000 ;
        RECT 116.490 165.650 117.300 165.920 ;
        RECT 116.490 165.380 117.030 165.650 ;
        RECT 116.760 165.110 117.030 165.380 ;
        RECT 118.110 165.110 118.920 165.920 ;
        RECT 119.730 165.650 120.540 165.920 ;
        RECT 120.000 165.380 120.540 165.650 ;
        RECT 120.000 165.110 120.270 165.380 ;
        RECT 116.760 164.840 117.300 165.110 ;
        RECT 117.840 164.840 119.190 165.110 ;
        RECT 119.730 164.840 120.270 165.110 ;
        RECT 116.760 164.570 118.380 164.840 ;
        RECT 118.650 164.570 120.000 164.840 ;
        RECT 117.300 164.300 118.110 164.570 ;
        RECT 118.920 164.300 120.000 164.570 ;
        RECT 117.570 163.760 119.460 164.300 ;
        RECT 115.950 163.490 116.760 163.760 ;
        RECT 117.570 163.490 117.840 163.760 ;
        RECT 118.110 163.490 118.380 163.760 ;
        RECT 118.650 163.490 118.920 163.760 ;
        RECT 119.190 163.490 119.460 163.760 ;
        RECT 120.270 163.490 121.080 163.760 ;
        RECT 115.680 162.950 117.030 163.490 ;
        RECT 120.000 162.950 121.350 163.490 ;
        RECT 115.950 162.680 117.570 162.950 ;
        RECT 119.460 162.680 121.080 162.950 ;
        RECT 116.760 162.410 117.840 162.680 ;
        RECT 119.190 162.410 120.270 162.680 ;
        RECT 114.890 162.135 115.840 162.410 ;
        RECT 117.300 162.140 118.380 162.410 ;
        RECT 118.650 162.140 119.730 162.410 ;
        RECT 121.340 162.265 122.340 162.410 ;
        RECT 47.950 161.220 49.200 161.620 ;
        RECT 49.370 161.260 52.880 161.800 ;
        RECT 110.265 161.585 115.840 162.135 ;
        RECT 117.840 161.600 119.190 162.140 ;
        RECT 121.340 161.715 123.765 162.265 ;
        RECT 114.890 161.510 115.840 161.585 ;
        RECT 117.300 161.330 118.380 161.600 ;
        RECT 118.650 161.330 119.730 161.600 ;
        RECT 121.340 161.510 122.340 161.715 ;
        RECT 47.950 161.070 48.450 161.220 ;
        RECT 49.910 160.990 52.340 161.260 ;
        RECT 115.950 161.060 117.840 161.330 ;
        RECT 119.190 161.060 121.350 161.330 ;
        RECT 50.180 160.720 52.340 160.990 ;
        RECT 115.680 160.790 117.300 161.060 ;
        RECT 119.730 160.790 121.350 161.060 ;
        RECT 115.680 160.520 116.760 160.790 ;
        RECT 120.270 160.520 121.350 160.790 ;
        RECT 115.680 160.250 116.490 160.520 ;
        RECT 120.540 160.250 121.350 160.520 ;
        RECT 115.950 159.980 116.220 160.250 ;
        RECT 117.570 159.980 117.840 160.250 ;
        RECT 118.110 159.980 118.380 160.250 ;
        RECT 118.650 159.980 118.920 160.250 ;
        RECT 119.190 159.980 119.460 160.250 ;
        RECT 120.810 159.980 121.080 160.250 ;
        RECT 117.570 159.440 119.460 159.980 ;
        RECT 117.300 159.170 118.110 159.440 ;
        RECT 118.920 159.170 120.000 159.440 ;
        RECT 116.760 158.900 118.380 159.170 ;
        RECT 118.650 158.900 120.000 159.170 ;
        RECT 116.760 158.630 117.300 158.900 ;
        RECT 117.840 158.630 119.190 158.900 ;
        RECT 119.730 158.630 120.270 158.900 ;
        RECT 116.760 158.360 117.030 158.630 ;
        RECT 116.490 158.090 117.030 158.360 ;
        RECT 116.490 157.820 117.300 158.090 ;
        RECT 118.110 157.820 118.920 158.630 ;
        RECT 120.000 158.360 120.270 158.630 ;
        RECT 120.000 158.090 120.540 158.360 ;
        RECT 119.730 157.820 120.540 158.090 ;
        RECT 116.490 156.740 120.540 157.820 ;
        RECT 26.120 146.940 28.280 147.210 ;
        RECT 23.890 146.690 24.290 146.790 ;
        RECT 23.890 146.240 24.890 146.690 ;
        RECT 25.850 146.670 28.280 146.940 ;
        RECT 25.310 146.130 28.820 146.670 ;
        RECT 25.040 145.050 29.090 146.130 ;
        RECT 25.040 144.780 25.850 145.050 ;
        RECT 25.040 144.510 25.580 144.780 ;
        RECT 25.310 144.240 25.580 144.510 ;
        RECT 26.660 144.240 27.470 145.050 ;
        RECT 28.280 144.780 29.090 145.050 ;
        RECT 28.550 144.510 29.090 144.780 ;
        RECT 28.550 144.240 28.820 144.510 ;
        RECT 25.310 143.970 25.850 144.240 ;
        RECT 26.390 143.970 27.740 144.240 ;
        RECT 28.280 143.970 28.820 144.240 ;
        RECT 25.310 143.700 26.930 143.970 ;
        RECT 27.200 143.700 28.550 143.970 ;
        RECT 25.850 143.430 26.660 143.700 ;
        RECT 27.470 143.430 28.550 143.700 ;
        RECT 26.120 142.890 28.010 143.430 ;
        RECT 24.500 142.620 25.310 142.890 ;
        RECT 26.120 142.620 26.390 142.890 ;
        RECT 26.660 142.620 26.930 142.890 ;
        RECT 27.200 142.620 27.470 142.890 ;
        RECT 27.740 142.620 28.010 142.890 ;
        RECT 28.820 142.620 29.630 142.890 ;
        RECT 24.230 142.080 25.580 142.620 ;
        RECT 28.550 142.080 29.900 142.620 ;
        RECT 24.500 141.810 26.120 142.080 ;
        RECT 28.010 141.810 29.630 142.080 ;
        RECT 25.310 141.540 26.390 141.810 ;
        RECT 27.740 141.540 28.820 141.810 ;
        RECT 30.880 141.540 31.380 155.600 ;
        RECT 33.510 155.420 34.460 155.600 ;
        RECT 36.460 155.510 37.810 156.050 ;
        RECT 39.960 155.630 43.710 156.130 ;
        RECT 115.340 156.160 116.590 156.560 ;
        RECT 116.760 156.200 120.270 156.740 ;
        RECT 115.340 156.010 115.840 156.160 ;
        RECT 117.300 155.930 119.730 156.200 ;
        RECT 117.570 155.660 119.730 155.930 ;
        RECT 35.920 155.240 37.000 155.510 ;
        RECT 37.270 155.240 38.350 155.510 ;
        RECT 39.960 155.420 40.960 155.630 ;
        RECT 34.570 154.970 36.460 155.240 ;
        RECT 37.810 154.970 39.970 155.240 ;
        RECT 34.300 154.700 35.920 154.970 ;
        RECT 38.350 154.700 39.970 154.970 ;
        RECT 34.300 154.430 35.380 154.700 ;
        RECT 38.890 154.430 39.970 154.700 ;
        RECT 34.300 154.160 35.110 154.430 ;
        RECT 39.160 154.160 39.970 154.430 ;
        RECT 34.570 153.890 34.840 154.160 ;
        RECT 36.190 153.890 36.460 154.160 ;
        RECT 36.730 153.890 37.000 154.160 ;
        RECT 37.270 153.890 37.540 154.160 ;
        RECT 37.810 153.890 38.080 154.160 ;
        RECT 39.430 153.890 39.700 154.160 ;
        RECT 36.190 153.350 38.080 153.890 ;
        RECT 35.920 153.080 36.730 153.350 ;
        RECT 37.540 153.080 38.620 153.350 ;
        RECT 35.380 152.810 37.000 153.080 ;
        RECT 37.270 152.810 38.620 153.080 ;
        RECT 35.380 152.540 35.920 152.810 ;
        RECT 36.460 152.540 37.810 152.810 ;
        RECT 38.350 152.540 38.890 152.810 ;
        RECT 35.380 152.270 35.650 152.540 ;
        RECT 35.110 152.000 35.650 152.270 ;
        RECT 35.110 151.730 35.920 152.000 ;
        RECT 36.730 151.730 37.540 152.540 ;
        RECT 38.620 152.270 38.890 152.540 ;
        RECT 38.620 152.000 39.160 152.270 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 38.350 151.730 39.160 152.000 ;
        RECT 35.110 150.650 39.160 151.730 ;
        RECT 33.960 150.070 35.210 150.470 ;
        RECT 35.380 150.110 38.890 150.650 ;
        RECT 33.960 149.920 34.460 150.070 ;
        RECT 35.920 149.840 38.350 150.110 ;
        RECT 36.190 149.570 38.350 149.840 ;
        RECT 68.170 149.600 91.570 152.200 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 123.215 149.205 123.765 161.715 ;
        RECT 129.740 154.700 131.900 154.970 ;
        RECT 127.510 154.450 127.910 154.550 ;
        RECT 127.510 154.000 128.510 154.450 ;
        RECT 129.470 154.430 131.900 154.700 ;
        RECT 128.930 153.890 132.440 154.430 ;
        RECT 128.660 152.810 132.710 153.890 ;
        RECT 128.660 152.540 129.470 152.810 ;
        RECT 128.660 152.270 129.200 152.540 ;
        RECT 128.930 152.000 129.200 152.270 ;
        RECT 130.280 152.000 131.090 152.810 ;
        RECT 131.900 152.540 132.710 152.810 ;
        RECT 132.170 152.270 132.710 152.540 ;
        RECT 132.170 152.000 132.440 152.270 ;
        RECT 128.930 151.730 129.470 152.000 ;
        RECT 130.010 151.730 131.360 152.000 ;
        RECT 131.900 151.730 132.440 152.000 ;
        RECT 128.930 151.460 130.550 151.730 ;
        RECT 130.820 151.460 132.170 151.730 ;
        RECT 129.470 151.190 130.280 151.460 ;
        RECT 131.090 151.190 132.170 151.460 ;
        RECT 129.740 150.650 131.630 151.190 ;
        RECT 128.120 150.380 128.930 150.650 ;
        RECT 129.740 150.380 130.010 150.650 ;
        RECT 130.280 150.380 130.550 150.650 ;
        RECT 130.820 150.380 131.090 150.650 ;
        RECT 131.360 150.380 131.630 150.650 ;
        RECT 132.440 150.380 133.250 150.650 ;
        RECT 127.850 149.840 129.200 150.380 ;
        RECT 132.170 149.840 133.520 150.380 ;
        RECT 128.120 149.570 129.740 149.840 ;
        RECT 131.630 149.570 133.250 149.840 ;
        RECT 128.930 149.300 130.010 149.570 ;
        RECT 131.360 149.300 132.440 149.570 ;
        RECT 127.060 149.205 128.010 149.300 ;
        RECT 123.215 148.655 128.010 149.205 ;
        RECT 129.470 149.030 130.550 149.300 ;
        RECT 130.820 149.030 131.900 149.300 ;
        RECT 133.510 149.075 134.510 149.300 ;
        RECT 127.060 148.400 128.010 148.655 ;
        RECT 130.010 148.490 131.360 149.030 ;
        RECT 133.510 148.525 135.725 149.075 ;
        RECT 129.470 148.220 130.550 148.490 ;
        RECT 130.820 148.220 131.900 148.490 ;
        RECT 133.510 148.400 134.510 148.525 ;
        RECT 128.120 147.950 130.010 148.220 ;
        RECT 131.360 147.950 133.520 148.220 ;
        RECT 127.850 147.680 129.470 147.950 ;
        RECT 131.900 147.680 133.520 147.950 ;
        RECT 127.850 147.410 128.930 147.680 ;
        RECT 132.440 147.410 133.520 147.680 ;
        RECT 127.850 147.140 128.660 147.410 ;
        RECT 132.710 147.140 133.520 147.410 ;
        RECT 128.120 146.870 128.390 147.140 ;
        RECT 129.740 146.870 130.010 147.140 ;
        RECT 130.280 146.870 130.550 147.140 ;
        RECT 130.820 146.870 131.090 147.140 ;
        RECT 131.360 146.870 131.630 147.140 ;
        RECT 132.980 146.870 133.250 147.140 ;
        RECT 129.740 146.330 131.630 146.870 ;
        RECT 129.470 146.060 130.280 146.330 ;
        RECT 131.090 146.060 132.170 146.330 ;
        RECT 128.930 145.790 130.550 146.060 ;
        RECT 130.820 145.790 132.170 146.060 ;
        RECT 128.930 145.520 129.470 145.790 ;
        RECT 130.010 145.520 131.360 145.790 ;
        RECT 131.900 145.520 132.440 145.790 ;
        RECT 128.930 145.250 129.200 145.520 ;
        RECT 128.660 144.980 129.200 145.250 ;
        RECT 128.660 144.710 129.470 144.980 ;
        RECT 130.280 144.710 131.090 145.520 ;
        RECT 132.170 145.250 132.440 145.520 ;
        RECT 132.170 144.980 132.710 145.250 ;
        RECT 131.900 144.710 132.710 144.980 ;
        RECT 23.440 141.300 24.390 141.540 ;
        RECT 17.400 140.800 24.390 141.300 ;
        RECT 25.850 141.270 26.930 141.540 ;
        RECT 27.200 141.270 28.280 141.540 ;
        RECT 17.400 124.190 17.900 140.800 ;
        RECT 23.440 140.640 24.390 140.800 ;
        RECT 26.390 140.730 27.740 141.270 ;
        RECT 29.890 140.850 31.380 141.540 ;
        RECT 25.850 140.460 26.930 140.730 ;
        RECT 27.200 140.460 28.280 140.730 ;
        RECT 29.890 140.640 30.890 140.850 ;
        RECT 24.500 140.190 26.390 140.460 ;
        RECT 27.740 140.190 29.900 140.460 ;
        RECT 24.230 139.920 25.850 140.190 ;
        RECT 28.280 139.920 29.900 140.190 ;
        RECT 24.230 139.650 25.310 139.920 ;
        RECT 28.820 139.650 29.900 139.920 ;
        RECT 24.230 139.380 25.040 139.650 ;
        RECT 29.090 139.380 29.900 139.650 ;
        RECT 24.500 139.110 24.770 139.380 ;
        RECT 26.120 139.110 26.390 139.380 ;
        RECT 26.660 139.110 26.930 139.380 ;
        RECT 27.200 139.110 27.470 139.380 ;
        RECT 27.740 139.110 28.010 139.380 ;
        RECT 29.360 139.110 29.630 139.380 ;
        RECT 26.120 138.570 28.010 139.110 ;
        RECT 25.850 138.300 26.660 138.570 ;
        RECT 27.470 138.300 28.550 138.570 ;
        RECT 25.310 138.030 26.930 138.300 ;
        RECT 27.200 138.030 28.550 138.300 ;
        RECT 25.310 137.760 25.850 138.030 ;
        RECT 26.390 137.760 27.740 138.030 ;
        RECT 28.280 137.760 28.820 138.030 ;
        RECT 25.310 137.490 25.580 137.760 ;
        RECT 25.040 137.220 25.580 137.490 ;
        RECT 25.040 136.950 25.850 137.220 ;
        RECT 26.660 136.950 27.470 137.760 ;
        RECT 28.550 137.490 28.820 137.760 ;
        RECT 28.550 137.220 29.090 137.490 ;
        RECT 28.280 136.950 29.090 137.220 ;
        RECT 25.040 135.870 29.090 136.950 ;
        RECT 23.890 135.290 25.140 135.690 ;
        RECT 25.310 135.330 28.820 135.870 ;
        RECT 23.890 135.140 24.390 135.290 ;
        RECT 25.850 135.060 28.280 135.330 ;
        RECT 26.120 134.790 28.280 135.060 ;
        RECT 60.370 134.000 99.370 144.400 ;
        RECT 128.660 143.630 132.710 144.710 ;
        RECT 127.510 143.050 128.760 143.450 ;
        RECT 128.930 143.090 132.440 143.630 ;
        RECT 127.510 142.900 128.010 143.050 ;
        RECT 129.470 142.820 131.900 143.090 ;
        RECT 129.740 142.550 131.900 142.820 ;
        RECT 135.175 142.355 135.725 148.525 ;
        RECT 135.175 141.805 143.285 142.355 ;
        RECT 137.430 138.590 139.590 138.860 ;
        RECT 137.430 138.320 139.860 138.590 ;
        RECT 141.420 138.340 141.820 138.440 ;
        RECT 136.890 137.780 140.400 138.320 ;
        RECT 140.820 137.890 141.820 138.340 ;
        RECT 136.620 136.700 140.670 137.780 ;
        RECT 136.620 136.430 137.430 136.700 ;
        RECT 136.620 136.160 137.160 136.430 ;
        RECT 136.890 135.890 137.160 136.160 ;
        RECT 138.240 135.890 139.050 136.700 ;
        RECT 139.860 136.430 140.670 136.700 ;
        RECT 140.130 136.160 140.670 136.430 ;
        RECT 140.130 135.890 140.400 136.160 ;
        RECT 136.890 135.620 137.430 135.890 ;
        RECT 137.970 135.620 139.320 135.890 ;
        RECT 139.860 135.620 140.400 135.890 ;
        RECT 137.160 135.350 138.510 135.620 ;
        RECT 138.780 135.350 140.400 135.620 ;
        RECT 137.160 135.080 138.240 135.350 ;
        RECT 139.050 135.080 139.860 135.350 ;
        RECT 137.700 134.540 139.590 135.080 ;
        RECT 136.080 134.270 136.890 134.540 ;
        RECT 137.700 134.270 137.970 134.540 ;
        RECT 138.240 134.270 138.510 134.540 ;
        RECT 138.780 134.270 139.050 134.540 ;
        RECT 139.320 134.270 139.590 134.540 ;
        RECT 140.400 134.270 141.210 134.540 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 20.780 129.850 22.940 130.120 ;
        RECT 20.780 129.580 23.210 129.850 ;
        RECT 24.770 129.600 25.170 129.700 ;
        RECT 20.240 129.040 23.750 129.580 ;
        RECT 24.170 129.150 25.170 129.600 ;
        RECT 19.970 127.960 24.020 129.040 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 19.970 127.690 20.780 127.960 ;
        RECT 19.970 127.420 20.510 127.690 ;
        RECT 20.240 127.150 20.510 127.420 ;
        RECT 21.590 127.150 22.400 127.960 ;
        RECT 23.210 127.690 24.020 127.960 ;
        RECT 23.480 127.420 24.020 127.690 ;
        RECT 23.480 127.150 23.750 127.420 ;
        RECT 20.240 126.880 20.780 127.150 ;
        RECT 21.320 126.880 22.670 127.150 ;
        RECT 23.210 126.880 23.750 127.150 ;
        RECT 20.510 126.610 21.860 126.880 ;
        RECT 22.130 126.610 23.750 126.880 ;
        RECT 20.510 126.340 21.590 126.610 ;
        RECT 22.400 126.340 23.210 126.610 ;
        RECT 21.050 125.800 22.940 126.340 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 135.810 133.730 137.160 134.270 ;
        RECT 140.130 133.730 141.480 134.270 ;
        RECT 136.080 133.460 137.700 133.730 ;
        RECT 139.590 133.460 141.210 133.730 ;
        RECT 136.890 133.190 137.970 133.460 ;
        RECT 139.320 133.190 140.400 133.460 ;
        RECT 134.820 132.990 135.820 133.190 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 134.120 132.490 135.820 132.990 ;
        RECT 137.430 132.920 138.510 133.190 ;
        RECT 138.780 132.920 139.860 133.190 ;
        RECT 141.320 133.115 142.270 133.190 ;
        RECT 142.735 133.115 143.285 141.805 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 19.430 125.530 20.240 125.800 ;
        RECT 21.050 125.530 21.320 125.800 ;
        RECT 21.590 125.530 21.860 125.800 ;
        RECT 22.130 125.530 22.400 125.800 ;
        RECT 22.670 125.530 22.940 125.800 ;
        RECT 23.750 125.530 24.560 125.800 ;
        RECT 19.160 124.990 20.510 125.530 ;
        RECT 23.480 124.990 24.830 125.530 ;
        RECT 19.430 124.720 21.050 124.990 ;
        RECT 22.940 124.720 24.560 124.990 ;
        RECT 20.240 124.450 21.320 124.720 ;
        RECT 22.670 124.450 23.750 124.720 ;
        RECT 18.170 124.190 19.170 124.450 ;
        RECT 17.400 123.690 19.170 124.190 ;
        RECT 20.780 124.180 21.860 124.450 ;
        RECT 22.130 124.180 23.210 124.450 ;
        RECT 24.670 124.290 25.620 124.450 ;
        RECT 18.170 123.550 19.170 123.690 ;
        RECT 21.320 123.640 22.670 124.180 ;
        RECT 24.670 123.790 26.800 124.290 ;
        RECT 20.780 123.370 21.860 123.640 ;
        RECT 22.130 123.370 23.210 123.640 ;
        RECT 24.670 123.550 25.620 123.790 ;
        RECT 19.160 123.100 21.320 123.370 ;
        RECT 22.670 123.100 24.560 123.370 ;
        RECT 19.160 122.830 20.780 123.100 ;
        RECT 23.210 122.830 24.830 123.100 ;
        RECT 19.160 122.560 20.240 122.830 ;
        RECT 23.750 122.560 24.830 122.830 ;
        RECT 19.160 122.290 19.970 122.560 ;
        RECT 24.020 122.290 24.830 122.560 ;
        RECT 19.430 122.020 19.700 122.290 ;
        RECT 21.050 122.020 21.320 122.290 ;
        RECT 21.590 122.020 21.860 122.290 ;
        RECT 22.130 122.020 22.400 122.290 ;
        RECT 22.670 122.020 22.940 122.290 ;
        RECT 24.290 122.020 24.560 122.290 ;
        RECT 21.050 121.480 22.940 122.020 ;
        RECT 20.510 121.210 21.590 121.480 ;
        RECT 22.400 121.210 23.210 121.480 ;
        RECT 20.510 120.940 21.860 121.210 ;
        RECT 22.130 120.940 23.750 121.210 ;
        RECT 20.240 120.670 20.780 120.940 ;
        RECT 21.320 120.670 22.670 120.940 ;
        RECT 23.210 120.670 23.750 120.940 ;
        RECT 20.240 120.400 20.510 120.670 ;
        RECT 19.970 120.130 20.510 120.400 ;
        RECT 19.970 119.860 20.780 120.130 ;
        RECT 21.590 119.860 22.400 120.670 ;
        RECT 23.480 120.400 23.750 120.670 ;
        RECT 23.480 120.130 24.020 120.400 ;
        RECT 23.210 119.860 24.020 120.130 ;
        RECT 19.970 118.780 24.020 119.860 ;
        RECT 20.240 118.240 23.750 118.780 ;
        RECT 20.780 117.970 23.210 118.240 ;
        RECT 23.920 118.200 25.170 118.600 ;
        RECT 24.670 118.050 25.170 118.200 ;
        RECT 20.780 117.700 22.940 117.970 ;
        RECT 7.470 112.910 9.070 114.410 ;
        RECT 20.850 111.970 23.010 112.240 ;
        RECT 18.620 111.720 19.020 111.820 ;
        RECT 18.620 111.270 19.620 111.720 ;
        RECT 20.580 111.700 23.010 111.970 ;
        RECT 20.040 111.160 23.550 111.700 ;
        RECT 19.770 110.080 23.820 111.160 ;
        RECT 19.770 109.810 20.580 110.080 ;
        RECT 19.770 109.540 20.310 109.810 ;
        RECT 20.040 109.270 20.310 109.540 ;
        RECT 21.390 109.270 22.200 110.080 ;
        RECT 23.010 109.810 23.820 110.080 ;
        RECT 23.280 109.540 23.820 109.810 ;
        RECT 23.280 109.270 23.550 109.540 ;
        RECT 20.040 109.000 20.580 109.270 ;
        RECT 21.120 109.000 22.470 109.270 ;
        RECT 23.010 109.000 23.550 109.270 ;
        RECT 20.040 108.730 21.660 109.000 ;
        RECT 21.930 108.730 23.280 109.000 ;
        RECT 20.580 108.460 21.390 108.730 ;
        RECT 22.200 108.460 23.280 108.730 ;
        RECT 20.850 107.920 22.740 108.460 ;
        RECT 19.230 107.650 20.040 107.920 ;
        RECT 20.850 107.650 21.120 107.920 ;
        RECT 21.390 107.650 21.660 107.920 ;
        RECT 21.930 107.650 22.200 107.920 ;
        RECT 22.470 107.650 22.740 107.920 ;
        RECT 23.550 107.650 24.360 107.920 ;
        RECT 18.960 107.110 20.310 107.650 ;
        RECT 23.280 107.110 24.630 107.650 ;
        RECT 19.230 106.840 20.850 107.110 ;
        RECT 22.740 106.840 24.360 107.110 ;
        RECT 20.040 106.570 21.120 106.840 ;
        RECT 22.470 106.570 23.550 106.840 ;
        RECT 18.170 106.360 19.120 106.570 ;
        RECT 17.240 105.860 19.120 106.360 ;
        RECT 20.580 106.300 21.660 106.570 ;
        RECT 21.930 106.300 23.010 106.570 ;
        RECT 24.620 106.370 25.620 106.570 ;
        RECT 26.300 106.370 26.800 123.790 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 30.710 114.330 31.810 115.530 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 134.120 115.250 134.620 132.490 ;
        RECT 134.820 132.290 135.820 132.490 ;
        RECT 137.970 132.380 139.320 132.920 ;
        RECT 141.320 132.565 143.285 133.115 ;
        RECT 137.430 132.110 138.510 132.380 ;
        RECT 138.780 132.110 139.860 132.380 ;
        RECT 141.320 132.290 142.270 132.565 ;
        RECT 135.810 131.840 137.970 132.110 ;
        RECT 139.320 131.840 141.210 132.110 ;
        RECT 135.810 131.570 137.430 131.840 ;
        RECT 139.860 131.570 141.480 131.840 ;
        RECT 135.810 131.300 136.890 131.570 ;
        RECT 140.400 131.300 141.480 131.570 ;
        RECT 135.810 131.030 136.620 131.300 ;
        RECT 140.670 131.030 141.480 131.300 ;
        RECT 136.080 130.760 136.350 131.030 ;
        RECT 137.700 130.760 137.970 131.030 ;
        RECT 138.240 130.760 138.510 131.030 ;
        RECT 138.780 130.760 139.050 131.030 ;
        RECT 139.320 130.760 139.590 131.030 ;
        RECT 140.940 130.760 141.210 131.030 ;
        RECT 137.700 130.220 139.590 130.760 ;
        RECT 137.160 129.950 138.240 130.220 ;
        RECT 139.050 129.950 139.860 130.220 ;
        RECT 137.160 129.680 138.510 129.950 ;
        RECT 138.780 129.680 140.400 129.950 ;
        RECT 136.890 129.410 137.430 129.680 ;
        RECT 137.970 129.410 139.320 129.680 ;
        RECT 139.860 129.410 140.400 129.680 ;
        RECT 136.890 129.140 137.160 129.410 ;
        RECT 136.620 128.870 137.160 129.140 ;
        RECT 136.620 128.600 137.430 128.870 ;
        RECT 138.240 128.600 139.050 129.410 ;
        RECT 140.130 129.140 140.400 129.410 ;
        RECT 140.130 128.870 140.670 129.140 ;
        RECT 139.860 128.600 140.670 128.870 ;
        RECT 136.620 127.520 140.670 128.600 ;
        RECT 136.890 126.980 140.400 127.520 ;
        RECT 137.430 126.710 139.860 126.980 ;
        RECT 140.570 126.940 141.820 127.340 ;
        RECT 141.320 126.790 141.820 126.940 ;
        RECT 137.430 126.440 139.590 126.710 ;
        RECT 140.170 120.910 142.330 121.180 ;
        RECT 137.940 120.660 138.340 120.760 ;
        RECT 137.940 120.210 138.940 120.660 ;
        RECT 139.900 120.640 142.330 120.910 ;
        RECT 139.360 120.100 142.870 120.640 ;
        RECT 139.090 119.020 143.140 120.100 ;
        RECT 139.090 118.750 139.900 119.020 ;
        RECT 139.090 118.480 139.630 118.750 ;
        RECT 139.360 118.210 139.630 118.480 ;
        RECT 140.710 118.210 141.520 119.020 ;
        RECT 142.330 118.750 143.140 119.020 ;
        RECT 142.600 118.480 143.140 118.750 ;
        RECT 142.600 118.210 142.870 118.480 ;
        RECT 139.360 117.940 139.900 118.210 ;
        RECT 140.440 117.940 141.790 118.210 ;
        RECT 142.330 117.940 142.870 118.210 ;
        RECT 139.360 117.670 140.980 117.940 ;
        RECT 141.250 117.670 142.600 117.940 ;
        RECT 139.900 117.400 140.710 117.670 ;
        RECT 141.520 117.400 142.600 117.670 ;
        RECT 140.170 116.860 142.060 117.400 ;
        RECT 138.550 116.590 139.360 116.860 ;
        RECT 140.170 116.590 140.440 116.860 ;
        RECT 140.710 116.590 140.980 116.860 ;
        RECT 141.250 116.590 141.520 116.860 ;
        RECT 141.790 116.590 142.060 116.860 ;
        RECT 142.870 116.590 143.680 116.860 ;
        RECT 138.280 116.050 139.630 116.590 ;
        RECT 142.600 116.050 143.950 116.590 ;
        RECT 138.550 115.780 140.170 116.050 ;
        RECT 142.060 115.780 143.680 116.050 ;
        RECT 139.360 115.510 140.440 115.780 ;
        RECT 141.790 115.510 142.870 115.780 ;
        RECT 137.490 115.250 138.440 115.510 ;
        RECT 134.120 114.750 138.440 115.250 ;
        RECT 139.900 115.240 140.980 115.510 ;
        RECT 141.250 115.240 142.330 115.510 ;
        RECT 143.940 115.300 144.940 115.510 ;
        RECT 137.490 114.610 138.440 114.750 ;
        RECT 140.440 114.700 141.790 115.240 ;
        RECT 143.940 114.800 145.740 115.300 ;
        RECT 139.900 114.430 140.980 114.700 ;
        RECT 141.250 114.430 142.330 114.700 ;
        RECT 143.940 114.610 144.940 114.800 ;
        RECT 138.550 114.160 140.440 114.430 ;
        RECT 141.790 114.160 143.950 114.430 ;
        RECT 138.280 113.890 139.900 114.160 ;
        RECT 142.330 113.890 143.950 114.160 ;
        RECT 138.280 113.620 139.360 113.890 ;
        RECT 142.870 113.620 143.950 113.890 ;
        RECT 138.280 113.350 139.090 113.620 ;
        RECT 143.140 113.350 143.950 113.620 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 138.550 113.080 138.820 113.350 ;
        RECT 140.170 113.080 140.440 113.350 ;
        RECT 140.710 113.080 140.980 113.350 ;
        RECT 141.250 113.080 141.520 113.350 ;
        RECT 141.790 113.080 142.060 113.350 ;
        RECT 143.410 113.080 143.680 113.350 ;
        RECT 140.170 112.540 142.060 113.080 ;
        RECT 139.900 112.270 140.710 112.540 ;
        RECT 141.520 112.270 142.600 112.540 ;
        RECT 139.360 112.000 140.980 112.270 ;
        RECT 141.250 112.000 142.600 112.270 ;
        RECT 139.360 111.730 139.900 112.000 ;
        RECT 140.440 111.730 141.790 112.000 ;
        RECT 142.330 111.730 142.870 112.000 ;
        RECT 139.360 111.460 139.630 111.730 ;
        RECT 139.090 111.190 139.630 111.460 ;
        RECT 139.090 110.920 139.900 111.190 ;
        RECT 140.710 110.920 141.520 111.730 ;
        RECT 142.600 111.460 142.870 111.730 ;
        RECT 142.600 111.190 143.140 111.460 ;
        RECT 142.330 110.920 143.140 111.190 ;
        RECT 17.240 89.210 17.740 105.860 ;
        RECT 18.170 105.670 19.120 105.860 ;
        RECT 21.120 105.760 22.470 106.300 ;
        RECT 24.620 105.870 26.800 106.370 ;
        RECT 20.580 105.490 21.660 105.760 ;
        RECT 21.930 105.490 23.010 105.760 ;
        RECT 24.620 105.670 25.620 105.870 ;
        RECT 19.230 105.220 21.120 105.490 ;
        RECT 22.470 105.220 24.630 105.490 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
        RECT 139.090 109.840 143.140 110.920 ;
        RECT 137.940 109.260 139.190 109.660 ;
        RECT 139.360 109.300 142.870 109.840 ;
        RECT 137.940 109.110 138.440 109.260 ;
        RECT 139.900 109.030 142.330 109.300 ;
        RECT 140.170 108.760 142.330 109.030 ;
        RECT 18.960 104.950 20.580 105.220 ;
        RECT 23.010 104.950 24.630 105.220 ;
        RECT 18.960 104.680 20.040 104.950 ;
        RECT 23.550 104.680 24.630 104.950 ;
        RECT 18.960 104.410 19.770 104.680 ;
        RECT 23.820 104.410 24.630 104.680 ;
        RECT 19.230 104.140 19.500 104.410 ;
        RECT 20.850 104.140 21.120 104.410 ;
        RECT 21.390 104.140 21.660 104.410 ;
        RECT 21.930 104.140 22.200 104.410 ;
        RECT 22.470 104.140 22.740 104.410 ;
        RECT 24.090 104.140 24.360 104.410 ;
        RECT 20.850 103.600 22.740 104.140 ;
        RECT 20.580 103.330 21.390 103.600 ;
        RECT 22.200 103.330 23.280 103.600 ;
        RECT 20.040 103.060 21.660 103.330 ;
        RECT 21.930 103.060 23.280 103.330 ;
        RECT 20.040 102.790 20.580 103.060 ;
        RECT 21.120 102.790 22.470 103.060 ;
        RECT 23.010 102.790 23.550 103.060 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 137.430 103.230 139.590 103.500 ;
        RECT 137.430 102.960 139.860 103.230 ;
        RECT 141.420 102.980 141.820 103.080 ;
        RECT 20.040 102.520 20.310 102.790 ;
        RECT 19.770 102.250 20.310 102.520 ;
        RECT 19.770 101.980 20.580 102.250 ;
        RECT 21.390 101.980 22.200 102.790 ;
        RECT 23.280 102.520 23.550 102.790 ;
        RECT 23.280 102.250 23.820 102.520 ;
        RECT 23.010 101.980 23.820 102.250 ;
        RECT 19.770 100.900 23.820 101.980 ;
        RECT 18.620 100.320 19.870 100.720 ;
        RECT 20.040 100.360 23.550 100.900 ;
        RECT 18.620 100.170 19.120 100.320 ;
        RECT 20.580 100.090 23.010 100.360 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 136.890 102.420 140.400 102.960 ;
        RECT 140.820 102.530 141.820 102.980 ;
        RECT 136.620 101.340 140.670 102.420 ;
        RECT 136.620 101.070 137.430 101.340 ;
        RECT 136.620 100.800 137.160 101.070 ;
        RECT 136.890 100.530 137.160 100.800 ;
        RECT 138.240 100.530 139.050 101.340 ;
        RECT 139.860 101.070 140.670 101.340 ;
        RECT 140.130 100.800 140.670 101.070 ;
        RECT 140.130 100.530 140.400 100.800 ;
        RECT 136.890 100.260 137.430 100.530 ;
        RECT 137.970 100.260 139.320 100.530 ;
        RECT 139.860 100.260 140.400 100.530 ;
        RECT 20.850 99.820 23.010 100.090 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
        RECT 137.160 99.990 138.510 100.260 ;
        RECT 138.780 99.990 140.400 100.260 ;
        RECT 137.160 99.720 138.240 99.990 ;
        RECT 139.050 99.720 139.860 99.990 ;
        RECT 137.700 99.180 139.590 99.720 ;
        RECT 136.080 98.910 136.890 99.180 ;
        RECT 137.700 98.910 137.970 99.180 ;
        RECT 138.240 98.910 138.510 99.180 ;
        RECT 138.780 98.910 139.050 99.180 ;
        RECT 139.320 98.910 139.590 99.180 ;
        RECT 140.400 98.910 141.210 99.180 ;
        RECT 135.810 98.370 137.160 98.910 ;
        RECT 140.130 98.370 141.480 98.910 ;
        RECT 136.080 98.100 137.700 98.370 ;
        RECT 139.590 98.100 141.210 98.370 ;
        RECT 136.890 97.830 137.970 98.100 ;
        RECT 139.320 97.830 140.400 98.100 ;
        RECT 26.050 94.880 28.210 95.150 ;
        RECT 26.050 94.610 28.480 94.880 ;
        RECT 30.040 94.630 30.440 94.730 ;
        RECT 25.510 94.070 29.020 94.610 ;
        RECT 29.440 94.180 30.440 94.630 ;
        RECT 25.240 92.990 29.290 94.070 ;
        RECT 25.240 92.720 26.050 92.990 ;
        RECT 25.240 92.450 25.780 92.720 ;
        RECT 25.510 92.180 25.780 92.450 ;
        RECT 26.860 92.180 27.670 92.990 ;
        RECT 28.480 92.720 29.290 92.990 ;
        RECT 28.750 92.450 29.290 92.720 ;
        RECT 28.750 92.180 29.020 92.450 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 134.820 97.560 135.820 97.830 ;
        RECT 137.430 97.560 138.510 97.830 ;
        RECT 138.780 97.560 139.860 97.830 ;
        RECT 141.320 97.670 142.270 97.830 ;
        RECT 145.240 97.670 145.740 114.800 ;
        RECT 134.700 96.930 135.820 97.560 ;
        RECT 137.970 97.020 139.320 97.560 ;
        RECT 141.320 97.170 145.740 97.670 ;
        RECT 25.510 91.910 26.050 92.180 ;
        RECT 26.590 91.910 27.940 92.180 ;
        RECT 28.480 91.910 29.020 92.180 ;
        RECT 25.780 91.640 27.130 91.910 ;
        RECT 27.400 91.640 29.020 91.910 ;
        RECT 25.780 91.370 26.860 91.640 ;
        RECT 27.670 91.370 28.480 91.640 ;
        RECT 26.320 90.830 28.210 91.370 ;
        RECT 24.700 90.560 25.510 90.830 ;
        RECT 26.320 90.560 26.590 90.830 ;
        RECT 26.860 90.560 27.130 90.830 ;
        RECT 27.400 90.560 27.670 90.830 ;
        RECT 27.940 90.560 28.210 90.830 ;
        RECT 29.020 90.560 29.830 90.830 ;
        RECT 24.430 90.020 25.780 90.560 ;
        RECT 28.750 90.020 30.100 90.560 ;
        RECT 24.700 89.750 26.320 90.020 ;
        RECT 28.210 89.750 29.830 90.020 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
        RECT 25.510 89.480 26.590 89.750 ;
        RECT 27.940 89.480 29.020 89.750 ;
        RECT 23.440 89.210 24.440 89.480 ;
        RECT 26.050 89.210 27.130 89.480 ;
        RECT 27.400 89.210 28.480 89.480 ;
        RECT 29.940 89.290 30.890 89.480 ;
        RECT 17.240 88.710 24.440 89.210 ;
        RECT 23.440 88.580 24.440 88.710 ;
        RECT 26.590 88.670 27.940 89.210 ;
        RECT 29.940 88.790 31.880 89.290 ;
        RECT 26.050 88.400 27.130 88.670 ;
        RECT 27.400 88.400 28.480 88.670 ;
        RECT 29.940 88.580 30.890 88.790 ;
        RECT 24.430 88.130 26.590 88.400 ;
        RECT 27.940 88.130 29.830 88.400 ;
        RECT 24.430 87.860 26.050 88.130 ;
        RECT 28.480 87.860 30.100 88.130 ;
        RECT 24.430 87.590 25.510 87.860 ;
        RECT 29.020 87.590 30.100 87.860 ;
        RECT 24.430 87.320 25.240 87.590 ;
        RECT 29.290 87.320 30.100 87.590 ;
        RECT 24.700 87.050 24.970 87.320 ;
        RECT 26.320 87.050 26.590 87.320 ;
        RECT 26.860 87.050 27.130 87.320 ;
        RECT 27.400 87.050 27.670 87.320 ;
        RECT 27.940 87.050 28.210 87.320 ;
        RECT 29.560 87.050 29.830 87.320 ;
        RECT 26.320 86.510 28.210 87.050 ;
        RECT 25.780 86.240 26.860 86.510 ;
        RECT 27.670 86.240 28.480 86.510 ;
        RECT 25.780 85.970 27.130 86.240 ;
        RECT 27.400 85.970 29.020 86.240 ;
        RECT 25.510 85.700 26.050 85.970 ;
        RECT 26.590 85.700 27.940 85.970 ;
        RECT 28.480 85.700 29.020 85.970 ;
        RECT 25.510 85.430 25.780 85.700 ;
        RECT 25.240 85.160 25.780 85.430 ;
        RECT 25.240 84.890 26.050 85.160 ;
        RECT 26.860 84.890 27.670 85.700 ;
        RECT 28.750 85.430 29.020 85.700 ;
        RECT 28.750 85.160 29.290 85.430 ;
        RECT 28.480 84.890 29.290 85.160 ;
        RECT 25.240 83.810 29.290 84.890 ;
        RECT 25.510 83.270 29.020 83.810 ;
        RECT 26.050 83.000 28.480 83.270 ;
        RECT 29.190 83.230 30.440 83.630 ;
        RECT 29.940 83.080 30.440 83.230 ;
        RECT 26.050 82.730 28.210 83.000 ;
        RECT 31.380 74.470 31.880 88.790 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 129.670 87.120 131.830 87.390 ;
        RECT 129.670 86.850 132.100 87.120 ;
        RECT 133.660 86.870 134.060 86.970 ;
        RECT 129.130 86.310 132.640 86.850 ;
        RECT 133.060 86.420 134.060 86.870 ;
        RECT 128.860 85.230 132.910 86.310 ;
        RECT 128.860 84.960 129.670 85.230 ;
        RECT 128.860 84.690 129.400 84.960 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
        RECT 129.130 84.420 129.400 84.690 ;
        RECT 130.480 84.420 131.290 85.230 ;
        RECT 132.100 84.960 132.910 85.230 ;
        RECT 132.370 84.690 132.910 84.960 ;
        RECT 132.370 84.420 132.640 84.690 ;
        RECT 129.130 84.150 129.670 84.420 ;
        RECT 130.210 84.150 131.560 84.420 ;
        RECT 132.100 84.150 132.640 84.420 ;
        RECT 129.400 83.880 130.750 84.150 ;
        RECT 131.020 83.880 132.640 84.150 ;
        RECT 129.400 83.610 130.480 83.880 ;
        RECT 131.290 83.610 132.100 83.880 ;
        RECT 129.940 83.070 131.830 83.610 ;
        RECT 128.320 82.800 129.130 83.070 ;
        RECT 129.940 82.800 130.210 83.070 ;
        RECT 130.480 82.800 130.750 83.070 ;
        RECT 131.020 82.800 131.290 83.070 ;
        RECT 131.560 82.800 131.830 83.070 ;
        RECT 132.640 82.800 133.450 83.070 ;
        RECT 128.050 82.260 129.400 82.800 ;
        RECT 132.370 82.260 133.720 82.800 ;
        RECT 36.120 79.880 38.280 80.150 ;
        RECT 36.120 79.610 38.550 79.880 ;
        RECT 40.010 79.650 40.510 79.800 ;
        RECT 35.580 79.070 39.090 79.610 ;
        RECT 39.260 79.250 40.510 79.650 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 128.320 81.990 129.940 82.260 ;
        RECT 131.830 81.990 133.450 82.260 ;
        RECT 129.130 81.720 130.210 81.990 ;
        RECT 131.560 81.720 132.640 81.990 ;
        RECT 127.060 81.580 128.060 81.720 ;
        RECT 123.970 81.080 128.060 81.580 ;
        RECT 129.670 81.450 130.750 81.720 ;
        RECT 131.020 81.450 132.100 81.720 ;
        RECT 133.560 81.550 134.510 81.720 ;
        RECT 134.700 81.550 135.200 96.930 ;
        RECT 137.430 96.750 138.510 97.020 ;
        RECT 138.780 96.750 139.860 97.020 ;
        RECT 141.320 96.930 142.270 97.170 ;
        RECT 135.810 96.480 137.970 96.750 ;
        RECT 139.320 96.480 141.210 96.750 ;
        RECT 135.810 96.210 137.430 96.480 ;
        RECT 139.860 96.210 141.480 96.480 ;
        RECT 135.810 95.940 136.890 96.210 ;
        RECT 140.400 95.940 141.480 96.210 ;
        RECT 135.810 95.670 136.620 95.940 ;
        RECT 140.670 95.670 141.480 95.940 ;
        RECT 136.080 95.400 136.350 95.670 ;
        RECT 137.700 95.400 137.970 95.670 ;
        RECT 138.240 95.400 138.510 95.670 ;
        RECT 138.780 95.400 139.050 95.670 ;
        RECT 139.320 95.400 139.590 95.670 ;
        RECT 140.940 95.400 141.210 95.670 ;
        RECT 137.700 94.860 139.590 95.400 ;
        RECT 137.160 94.590 138.240 94.860 ;
        RECT 139.050 94.590 139.860 94.860 ;
        RECT 137.160 94.320 138.510 94.590 ;
        RECT 138.780 94.320 140.400 94.590 ;
        RECT 136.890 94.050 137.430 94.320 ;
        RECT 137.970 94.050 139.320 94.320 ;
        RECT 139.860 94.050 140.400 94.320 ;
        RECT 136.890 93.780 137.160 94.050 ;
        RECT 136.620 93.510 137.160 93.780 ;
        RECT 136.620 93.240 137.430 93.510 ;
        RECT 138.240 93.240 139.050 94.050 ;
        RECT 140.130 93.780 140.400 94.050 ;
        RECT 140.130 93.510 140.670 93.780 ;
        RECT 139.860 93.240 140.670 93.510 ;
        RECT 136.620 92.160 140.670 93.240 ;
        RECT 136.890 91.620 140.400 92.160 ;
        RECT 137.430 91.350 139.860 91.620 ;
        RECT 140.570 91.580 141.820 91.980 ;
        RECT 141.320 91.430 141.820 91.580 ;
        RECT 137.430 91.080 139.590 91.350 ;
        RECT 35.310 77.990 39.360 79.070 ;
        RECT 35.310 77.720 36.120 77.990 ;
        RECT 35.310 77.450 35.850 77.720 ;
        RECT 35.580 77.180 35.850 77.450 ;
        RECT 36.930 77.180 37.740 77.990 ;
        RECT 38.550 77.720 39.360 77.990 ;
        RECT 38.820 77.450 39.360 77.720 ;
        RECT 38.820 77.180 39.090 77.450 ;
        RECT 35.580 76.910 36.120 77.180 ;
        RECT 36.660 76.910 38.010 77.180 ;
        RECT 38.550 76.910 39.090 77.180 ;
        RECT 35.850 76.640 37.200 76.910 ;
        RECT 37.470 76.640 39.090 76.910 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
        RECT 35.850 76.370 36.930 76.640 ;
        RECT 37.740 76.370 38.550 76.640 ;
        RECT 36.390 75.830 38.280 76.370 ;
        RECT 34.770 75.560 35.040 75.830 ;
        RECT 36.390 75.560 36.660 75.830 ;
        RECT 36.930 75.560 37.200 75.830 ;
        RECT 37.470 75.560 37.740 75.830 ;
        RECT 38.010 75.560 38.280 75.830 ;
        RECT 39.630 75.560 39.900 75.830 ;
        RECT 34.500 75.290 35.310 75.560 ;
        RECT 39.360 75.290 40.170 75.560 ;
        RECT 34.500 75.020 35.580 75.290 ;
        RECT 39.090 75.020 40.170 75.290 ;
        RECT 34.500 74.750 36.120 75.020 ;
        RECT 38.550 74.750 40.170 75.020 ;
        RECT 34.500 74.480 36.660 74.750 ;
        RECT 38.010 74.480 39.900 74.750 ;
        RECT 31.380 74.300 33.950 74.470 ;
        RECT 31.380 73.970 34.510 74.300 ;
        RECT 36.120 74.210 37.200 74.480 ;
        RECT 37.470 74.210 38.550 74.480 ;
        RECT 40.460 74.300 43.980 74.520 ;
        RECT 33.510 73.400 34.510 73.970 ;
        RECT 36.660 73.670 38.010 74.210 ;
        RECT 40.010 74.020 43.980 74.300 ;
        RECT 36.120 73.400 37.200 73.670 ;
        RECT 37.470 73.400 38.550 73.670 ;
        RECT 40.010 73.400 40.960 74.020 ;
        RECT 35.580 73.130 36.660 73.400 ;
        RECT 38.010 73.130 39.090 73.400 ;
        RECT 34.770 72.860 36.390 73.130 ;
        RECT 38.280 72.860 39.900 73.130 ;
        RECT 34.500 72.320 35.850 72.860 ;
        RECT 38.820 72.320 40.170 72.860 ;
        RECT 34.770 72.050 35.580 72.320 ;
        RECT 36.390 72.050 36.660 72.320 ;
        RECT 36.930 72.050 37.200 72.320 ;
        RECT 37.470 72.050 37.740 72.320 ;
        RECT 38.010 72.050 38.280 72.320 ;
        RECT 39.090 72.050 39.900 72.320 ;
        RECT 36.390 71.510 38.280 72.050 ;
        RECT 35.850 71.240 36.930 71.510 ;
        RECT 37.740 71.240 38.550 71.510 ;
        RECT 35.850 70.970 37.200 71.240 ;
        RECT 37.470 70.970 39.090 71.240 ;
        RECT 35.580 70.700 36.120 70.970 ;
        RECT 36.660 70.700 38.010 70.970 ;
        RECT 38.550 70.700 39.090 70.970 ;
        RECT 35.580 70.430 35.850 70.700 ;
        RECT 35.310 70.160 35.850 70.430 ;
        RECT 35.310 69.890 36.120 70.160 ;
        RECT 36.930 69.890 37.740 70.700 ;
        RECT 38.820 70.430 39.090 70.700 ;
        RECT 38.820 70.160 39.360 70.430 ;
        RECT 38.550 69.890 39.360 70.160 ;
        RECT 35.310 68.810 39.360 69.890 ;
        RECT 35.580 68.270 39.090 68.810 ;
        RECT 36.120 68.000 38.550 68.270 ;
        RECT 39.510 68.250 40.510 68.700 ;
        RECT 40.110 68.150 40.510 68.250 ;
        RECT 36.120 67.730 38.280 68.000 ;
        RECT 43.480 63.340 43.980 74.020 ;
        RECT 117.500 73.790 119.660 74.060 ;
        RECT 117.500 73.520 119.930 73.790 ;
        RECT 121.390 73.560 121.890 73.710 ;
        RECT 116.960 72.980 120.470 73.520 ;
        RECT 120.640 73.160 121.890 73.560 ;
        RECT 116.690 71.900 120.740 72.980 ;
        RECT 116.690 71.630 117.500 71.900 ;
        RECT 116.690 71.360 117.230 71.630 ;
        RECT 116.960 71.090 117.230 71.360 ;
        RECT 118.310 71.090 119.120 71.900 ;
        RECT 119.930 71.630 120.740 71.900 ;
        RECT 120.200 71.360 120.740 71.630 ;
        RECT 120.200 71.090 120.470 71.360 ;
        RECT 116.960 70.820 117.500 71.090 ;
        RECT 118.040 70.820 119.390 71.090 ;
        RECT 119.930 70.820 120.470 71.090 ;
        RECT 117.230 70.550 118.580 70.820 ;
        RECT 118.850 70.550 120.470 70.820 ;
        RECT 117.230 70.280 118.310 70.550 ;
        RECT 119.120 70.280 119.930 70.550 ;
        RECT 117.770 69.740 119.660 70.280 ;
        RECT 116.150 69.470 116.420 69.740 ;
        RECT 117.770 69.470 118.040 69.740 ;
        RECT 118.310 69.470 118.580 69.740 ;
        RECT 118.850 69.470 119.120 69.740 ;
        RECT 119.390 69.470 119.660 69.740 ;
        RECT 121.010 69.470 121.280 69.740 ;
        RECT 115.880 69.200 116.690 69.470 ;
        RECT 120.740 69.200 121.550 69.470 ;
        RECT 50.100 68.730 52.260 69.000 ;
        RECT 115.880 68.930 116.960 69.200 ;
        RECT 120.470 68.930 121.550 69.200 ;
        RECT 50.100 68.460 52.530 68.730 ;
        RECT 115.880 68.660 117.500 68.930 ;
        RECT 119.930 68.660 121.550 68.930 ;
        RECT 53.990 68.500 54.490 68.650 ;
        RECT 49.560 67.920 53.070 68.460 ;
        RECT 53.240 68.100 54.490 68.500 ;
        RECT 115.880 68.390 118.040 68.660 ;
        RECT 119.390 68.390 121.280 68.660 ;
        RECT 123.970 68.390 124.470 81.080 ;
        RECT 127.060 80.820 128.060 81.080 ;
        RECT 130.210 80.910 131.560 81.450 ;
        RECT 133.560 81.050 135.200 81.550 ;
        RECT 129.670 80.640 130.750 80.910 ;
        RECT 131.020 80.640 132.100 80.910 ;
        RECT 133.560 80.820 134.510 81.050 ;
        RECT 128.050 80.370 130.210 80.640 ;
        RECT 131.560 80.370 133.450 80.640 ;
        RECT 128.050 80.100 129.670 80.370 ;
        RECT 132.100 80.100 133.720 80.370 ;
        RECT 128.050 79.830 129.130 80.100 ;
        RECT 132.640 79.830 133.720 80.100 ;
        RECT 128.050 79.560 128.860 79.830 ;
        RECT 132.910 79.560 133.720 79.830 ;
        RECT 128.320 79.290 128.590 79.560 ;
        RECT 129.940 79.290 130.210 79.560 ;
        RECT 130.480 79.290 130.750 79.560 ;
        RECT 131.020 79.290 131.290 79.560 ;
        RECT 131.560 79.290 131.830 79.560 ;
        RECT 133.180 79.290 133.450 79.560 ;
        RECT 129.940 78.750 131.830 79.290 ;
        RECT 129.400 78.480 130.480 78.750 ;
        RECT 131.290 78.480 132.100 78.750 ;
        RECT 129.400 78.210 130.750 78.480 ;
        RECT 131.020 78.210 132.640 78.480 ;
        RECT 129.130 77.940 129.670 78.210 ;
        RECT 130.210 77.940 131.560 78.210 ;
        RECT 132.100 77.940 132.640 78.210 ;
        RECT 129.130 77.670 129.400 77.940 ;
        RECT 128.860 77.400 129.400 77.670 ;
        RECT 128.860 77.130 129.670 77.400 ;
        RECT 130.480 77.130 131.290 77.940 ;
        RECT 132.370 77.670 132.640 77.940 ;
        RECT 132.370 77.400 132.910 77.670 ;
        RECT 132.100 77.130 132.910 77.400 ;
        RECT 128.860 76.050 132.910 77.130 ;
        RECT 129.130 75.510 132.640 76.050 ;
        RECT 129.670 75.240 132.100 75.510 ;
        RECT 132.810 75.470 134.060 75.870 ;
        RECT 133.560 75.320 134.060 75.470 ;
        RECT 129.670 74.970 131.830 75.240 ;
        RECT 109.160 68.210 115.260 68.340 ;
        RECT 49.290 66.840 53.340 67.920 ;
        RECT 49.290 66.570 50.100 66.840 ;
        RECT 49.290 66.300 49.830 66.570 ;
        RECT 49.560 66.030 49.830 66.300 ;
        RECT 50.910 66.030 51.720 66.840 ;
        RECT 52.530 66.570 53.340 66.840 ;
        RECT 52.800 66.300 53.340 66.570 ;
        RECT 109.160 67.840 115.890 68.210 ;
        RECT 117.500 68.120 118.580 68.390 ;
        RECT 118.850 68.120 119.930 68.390 ;
        RECT 121.840 68.210 124.470 68.390 ;
        RECT 52.800 66.030 53.070 66.300 ;
        RECT 49.560 65.760 50.100 66.030 ;
        RECT 50.640 65.760 51.990 66.030 ;
        RECT 52.530 65.760 53.070 66.030 ;
        RECT 49.830 65.490 51.180 65.760 ;
        RECT 51.450 65.490 53.070 65.760 ;
        RECT 49.830 65.220 50.910 65.490 ;
        RECT 51.720 65.220 52.530 65.490 ;
        RECT 50.370 64.680 52.260 65.220 ;
        RECT 102.020 64.840 104.180 65.110 ;
        RECT 48.750 64.410 49.020 64.680 ;
        RECT 50.370 64.410 50.640 64.680 ;
        RECT 50.910 64.410 51.180 64.680 ;
        RECT 51.450 64.410 51.720 64.680 ;
        RECT 51.990 64.410 52.260 64.680 ;
        RECT 53.610 64.410 53.880 64.680 ;
        RECT 102.020 64.570 104.450 64.840 ;
        RECT 105.910 64.610 106.410 64.760 ;
        RECT 48.480 64.140 49.290 64.410 ;
        RECT 53.340 64.140 54.150 64.410 ;
        RECT 48.480 63.870 49.560 64.140 ;
        RECT 53.070 63.870 54.150 64.140 ;
        RECT 101.480 64.030 104.990 64.570 ;
        RECT 105.160 64.210 106.410 64.610 ;
        RECT 48.480 63.600 50.100 63.870 ;
        RECT 52.530 63.600 54.150 63.870 ;
        RECT 43.480 63.150 47.690 63.340 ;
        RECT 48.480 63.330 50.640 63.600 ;
        RECT 51.990 63.330 53.880 63.600 ;
        RECT 43.480 62.840 48.490 63.150 ;
        RECT 50.100 63.060 51.180 63.330 ;
        RECT 51.450 63.060 52.530 63.330 ;
        RECT 54.440 63.150 56.740 63.440 ;
        RECT 47.490 62.250 48.490 62.840 ;
        RECT 50.640 62.520 51.990 63.060 ;
        RECT 53.990 62.940 56.740 63.150 ;
        RECT 50.100 62.250 51.180 62.520 ;
        RECT 51.450 62.250 52.530 62.520 ;
        RECT 53.990 62.250 54.940 62.940 ;
        RECT 49.560 61.980 50.640 62.250 ;
        RECT 51.990 61.980 53.070 62.250 ;
        RECT 48.750 61.710 50.370 61.980 ;
        RECT 52.260 61.710 53.880 61.980 ;
        RECT 48.480 61.170 49.830 61.710 ;
        RECT 52.800 61.170 54.150 61.710 ;
        RECT 48.750 60.900 49.560 61.170 ;
        RECT 50.370 60.900 50.640 61.170 ;
        RECT 50.910 60.900 51.180 61.170 ;
        RECT 51.450 60.900 51.720 61.170 ;
        RECT 51.990 60.900 52.260 61.170 ;
        RECT 53.070 60.900 53.880 61.170 ;
        RECT 50.370 60.360 52.260 60.900 ;
        RECT 49.830 60.090 50.910 60.360 ;
        RECT 51.720 60.090 52.530 60.360 ;
        RECT 49.830 59.820 51.180 60.090 ;
        RECT 51.450 59.820 53.070 60.090 ;
        RECT 49.560 59.550 50.100 59.820 ;
        RECT 50.640 59.550 51.990 59.820 ;
        RECT 52.530 59.550 53.070 59.820 ;
        RECT 49.560 59.280 49.830 59.550 ;
        RECT 49.290 59.010 49.830 59.280 ;
        RECT 49.290 58.740 50.100 59.010 ;
        RECT 50.910 58.740 51.720 59.550 ;
        RECT 52.800 59.280 53.070 59.550 ;
        RECT 52.800 59.010 53.340 59.280 ;
        RECT 52.530 58.740 53.340 59.010 ;
        RECT 49.290 57.660 53.340 58.740 ;
        RECT 49.560 57.120 53.070 57.660 ;
        RECT 50.100 56.850 52.530 57.120 ;
        RECT 53.490 57.100 54.490 57.550 ;
        RECT 54.090 57.000 54.490 57.100 ;
        RECT 56.240 56.910 56.740 62.940 ;
        RECT 101.210 62.950 105.260 64.030 ;
        RECT 101.210 62.680 102.020 62.950 ;
        RECT 66.750 62.200 68.910 62.470 ;
        RECT 101.210 62.410 101.750 62.680 ;
        RECT 66.750 61.930 69.180 62.200 ;
        RECT 101.480 62.140 101.750 62.410 ;
        RECT 102.830 62.140 103.640 62.950 ;
        RECT 104.450 62.680 105.260 62.950 ;
        RECT 104.720 62.410 105.260 62.680 ;
        RECT 104.720 62.140 104.990 62.410 ;
        RECT 70.640 61.970 71.140 62.120 ;
        RECT 66.210 61.390 69.720 61.930 ;
        RECT 69.890 61.570 71.140 61.970 ;
        RECT 101.480 61.870 102.020 62.140 ;
        RECT 102.560 61.870 103.910 62.140 ;
        RECT 104.450 61.870 104.990 62.140 ;
        RECT 101.750 61.600 103.100 61.870 ;
        RECT 103.370 61.600 104.990 61.870 ;
        RECT 65.940 60.310 69.990 61.390 ;
        RECT 101.750 61.330 102.830 61.600 ;
        RECT 103.640 61.330 104.450 61.600 ;
        RECT 84.580 60.860 86.740 61.130 ;
        RECT 84.580 60.590 87.010 60.860 ;
        RECT 102.290 60.790 104.180 61.330 ;
        RECT 88.470 60.630 88.970 60.780 ;
        RECT 65.940 60.040 66.750 60.310 ;
        RECT 65.940 59.770 66.480 60.040 ;
        RECT 66.210 59.500 66.480 59.770 ;
        RECT 67.560 59.500 68.370 60.310 ;
        RECT 69.180 60.040 69.990 60.310 ;
        RECT 84.040 60.050 87.550 60.590 ;
        RECT 87.720 60.230 88.970 60.630 ;
        RECT 100.670 60.520 100.940 60.790 ;
        RECT 102.290 60.520 102.560 60.790 ;
        RECT 102.830 60.520 103.100 60.790 ;
        RECT 103.370 60.520 103.640 60.790 ;
        RECT 103.910 60.520 104.180 60.790 ;
        RECT 105.530 60.520 105.800 60.790 ;
        RECT 100.400 60.250 101.210 60.520 ;
        RECT 105.260 60.250 106.070 60.520 ;
        RECT 69.450 59.770 69.990 60.040 ;
        RECT 69.450 59.500 69.720 59.770 ;
        RECT 66.210 59.230 66.750 59.500 ;
        RECT 67.290 59.230 68.640 59.500 ;
        RECT 69.180 59.230 69.720 59.500 ;
        RECT 66.480 58.960 67.830 59.230 ;
        RECT 68.100 58.960 69.720 59.230 ;
        RECT 83.770 58.970 87.820 60.050 ;
        RECT 100.400 59.980 101.480 60.250 ;
        RECT 104.990 59.980 106.070 60.250 ;
        RECT 100.400 59.710 102.020 59.980 ;
        RECT 104.450 59.710 106.070 59.980 ;
        RECT 66.480 58.690 67.560 58.960 ;
        RECT 68.370 58.690 69.180 58.960 ;
        RECT 83.770 58.700 84.580 58.970 ;
        RECT 67.020 58.150 68.910 58.690 ;
        RECT 83.770 58.430 84.310 58.700 ;
        RECT 84.040 58.160 84.310 58.430 ;
        RECT 85.390 58.160 86.200 58.970 ;
        RECT 87.010 58.700 87.820 58.970 ;
        RECT 87.280 58.430 87.820 58.700 ;
        RECT 92.210 59.260 99.720 59.520 ;
        RECT 100.400 59.440 102.560 59.710 ;
        RECT 103.910 59.440 105.800 59.710 ;
        RECT 109.160 59.440 109.660 67.840 ;
        RECT 114.890 67.310 115.890 67.840 ;
        RECT 118.040 67.580 119.390 68.120 ;
        RECT 121.390 67.890 124.470 68.210 ;
        RECT 117.500 67.310 118.580 67.580 ;
        RECT 118.850 67.310 119.930 67.580 ;
        RECT 121.390 67.310 122.340 67.890 ;
        RECT 116.960 67.040 118.040 67.310 ;
        RECT 119.390 67.040 120.470 67.310 ;
        RECT 116.150 66.770 117.770 67.040 ;
        RECT 119.660 66.770 121.280 67.040 ;
        RECT 115.880 66.230 117.230 66.770 ;
        RECT 120.200 66.230 121.550 66.770 ;
        RECT 116.150 65.960 116.960 66.230 ;
        RECT 117.770 65.960 118.040 66.230 ;
        RECT 118.310 65.960 118.580 66.230 ;
        RECT 118.850 65.960 119.120 66.230 ;
        RECT 119.390 65.960 119.660 66.230 ;
        RECT 120.470 65.960 121.280 66.230 ;
        RECT 117.770 65.420 119.660 65.960 ;
        RECT 117.230 65.150 118.310 65.420 ;
        RECT 119.120 65.150 119.930 65.420 ;
        RECT 117.230 64.880 118.580 65.150 ;
        RECT 118.850 64.880 120.470 65.150 ;
        RECT 116.960 64.610 117.500 64.880 ;
        RECT 118.040 64.610 119.390 64.880 ;
        RECT 119.930 64.610 120.470 64.880 ;
        RECT 116.960 64.340 117.230 64.610 ;
        RECT 116.690 64.070 117.230 64.340 ;
        RECT 116.690 63.800 117.500 64.070 ;
        RECT 118.310 63.800 119.120 64.610 ;
        RECT 120.200 64.340 120.470 64.610 ;
        RECT 120.200 64.070 120.740 64.340 ;
        RECT 119.930 63.800 120.740 64.070 ;
        RECT 116.690 62.720 120.740 63.800 ;
        RECT 116.960 62.180 120.470 62.720 ;
        RECT 117.500 61.910 119.930 62.180 ;
        RECT 120.890 62.160 121.890 62.610 ;
        RECT 121.490 62.060 121.890 62.160 ;
        RECT 117.500 61.640 119.660 61.910 ;
        RECT 92.210 59.020 100.410 59.260 ;
        RECT 102.020 59.170 103.100 59.440 ;
        RECT 103.370 59.170 104.450 59.440 ;
        RECT 106.360 59.260 109.660 59.440 ;
        RECT 87.280 58.160 87.550 58.430 ;
        RECT 65.400 57.880 65.670 58.150 ;
        RECT 67.020 57.880 67.290 58.150 ;
        RECT 67.560 57.880 67.830 58.150 ;
        RECT 68.100 57.880 68.370 58.150 ;
        RECT 68.640 57.880 68.910 58.150 ;
        RECT 70.260 57.880 70.530 58.150 ;
        RECT 84.040 57.890 84.580 58.160 ;
        RECT 85.120 57.890 86.470 58.160 ;
        RECT 87.010 57.890 87.550 58.160 ;
        RECT 65.130 57.610 65.940 57.880 ;
        RECT 69.990 57.610 70.800 57.880 ;
        RECT 65.130 57.340 66.210 57.610 ;
        RECT 69.720 57.340 70.800 57.610 ;
        RECT 84.310 57.620 85.660 57.890 ;
        RECT 85.930 57.620 87.550 57.890 ;
        RECT 84.310 57.350 85.390 57.620 ;
        RECT 86.200 57.350 87.010 57.620 ;
        RECT 65.130 57.070 66.750 57.340 ;
        RECT 69.180 57.070 70.800 57.340 ;
        RECT 50.100 56.580 52.260 56.850 ;
        RECT 56.240 56.620 64.470 56.910 ;
        RECT 65.130 56.800 67.290 57.070 ;
        RECT 68.640 56.800 70.530 57.070 ;
        RECT 56.240 56.410 65.140 56.620 ;
        RECT 66.750 56.530 67.830 56.800 ;
        RECT 68.100 56.530 69.180 56.800 ;
        RECT 71.090 56.620 76.900 56.820 ;
        RECT 84.850 56.810 86.740 57.350 ;
        RECT 64.140 55.720 65.140 56.410 ;
        RECT 67.290 55.990 68.640 56.530 ;
        RECT 70.640 56.320 76.900 56.620 ;
        RECT 83.230 56.540 83.500 56.810 ;
        RECT 84.850 56.540 85.120 56.810 ;
        RECT 85.390 56.540 85.660 56.810 ;
        RECT 85.930 56.540 86.200 56.810 ;
        RECT 86.470 56.540 86.740 56.810 ;
        RECT 88.090 56.540 88.360 56.810 ;
        RECT 66.750 55.720 67.830 55.990 ;
        RECT 68.100 55.720 69.180 55.990 ;
        RECT 70.640 55.720 71.590 56.320 ;
        RECT 66.210 55.450 67.290 55.720 ;
        RECT 68.640 55.450 69.720 55.720 ;
        RECT 76.400 55.460 76.900 56.320 ;
        RECT 82.960 56.270 83.770 56.540 ;
        RECT 87.820 56.270 88.630 56.540 ;
        RECT 82.960 56.000 84.040 56.270 ;
        RECT 87.550 56.000 88.630 56.270 ;
        RECT 82.960 55.730 84.580 56.000 ;
        RECT 87.010 55.730 88.630 56.000 ;
        RECT 82.960 55.460 85.120 55.730 ;
        RECT 86.470 55.460 88.360 55.730 ;
        RECT 65.400 55.180 67.020 55.450 ;
        RECT 68.910 55.180 70.530 55.450 ;
        RECT 76.400 55.280 82.320 55.460 ;
        RECT 65.130 54.640 66.480 55.180 ;
        RECT 69.450 54.640 70.800 55.180 ;
        RECT 76.400 54.960 82.970 55.280 ;
        RECT 84.580 55.190 85.660 55.460 ;
        RECT 85.930 55.190 87.010 55.460 ;
        RECT 92.210 55.440 92.710 59.020 ;
        RECT 99.410 58.360 100.410 59.020 ;
        RECT 102.560 58.630 103.910 59.170 ;
        RECT 105.910 58.940 109.660 59.260 ;
        RECT 102.020 58.360 103.100 58.630 ;
        RECT 103.370 58.360 104.450 58.630 ;
        RECT 105.910 58.360 106.860 58.940 ;
        RECT 101.480 58.090 102.560 58.360 ;
        RECT 103.910 58.090 104.990 58.360 ;
        RECT 100.670 57.820 102.290 58.090 ;
        RECT 104.180 57.820 105.800 58.090 ;
        RECT 100.400 57.280 101.750 57.820 ;
        RECT 104.720 57.280 106.070 57.820 ;
        RECT 100.670 57.010 101.480 57.280 ;
        RECT 102.290 57.010 102.560 57.280 ;
        RECT 102.830 57.010 103.100 57.280 ;
        RECT 103.370 57.010 103.640 57.280 ;
        RECT 103.910 57.010 104.180 57.280 ;
        RECT 104.990 57.010 105.800 57.280 ;
        RECT 102.290 56.470 104.180 57.010 ;
        RECT 101.750 56.200 102.830 56.470 ;
        RECT 103.640 56.200 104.450 56.470 ;
        RECT 101.750 55.930 103.100 56.200 ;
        RECT 103.370 55.930 104.990 56.200 ;
        RECT 88.920 55.280 92.710 55.440 ;
        RECT 101.480 55.660 102.020 55.930 ;
        RECT 102.560 55.660 103.910 55.930 ;
        RECT 104.450 55.660 104.990 55.930 ;
        RECT 101.480 55.390 101.750 55.660 ;
        RECT 65.400 54.370 66.210 54.640 ;
        RECT 67.020 54.370 67.290 54.640 ;
        RECT 67.560 54.370 67.830 54.640 ;
        RECT 68.100 54.370 68.370 54.640 ;
        RECT 68.640 54.370 68.910 54.640 ;
        RECT 69.720 54.370 70.530 54.640 ;
        RECT 81.970 54.380 82.970 54.960 ;
        RECT 85.120 54.650 86.470 55.190 ;
        RECT 88.470 54.940 92.710 55.280 ;
        RECT 101.210 55.120 101.750 55.390 ;
        RECT 84.580 54.380 85.660 54.650 ;
        RECT 85.930 54.380 87.010 54.650 ;
        RECT 88.470 54.380 89.420 54.940 ;
        RECT 101.210 54.850 102.020 55.120 ;
        RECT 102.830 54.850 103.640 55.660 ;
        RECT 104.720 55.390 104.990 55.660 ;
        RECT 104.720 55.120 105.260 55.390 ;
        RECT 104.450 54.850 105.260 55.120 ;
        RECT 67.020 53.830 68.910 54.370 ;
        RECT 84.040 54.110 85.120 54.380 ;
        RECT 86.470 54.110 87.550 54.380 ;
        RECT 83.230 53.840 84.850 54.110 ;
        RECT 86.740 53.840 88.360 54.110 ;
        RECT 66.480 53.560 67.560 53.830 ;
        RECT 68.370 53.560 69.180 53.830 ;
        RECT 66.480 53.290 67.830 53.560 ;
        RECT 68.100 53.290 69.720 53.560 ;
        RECT 82.960 53.300 84.310 53.840 ;
        RECT 87.280 53.300 88.630 53.840 ;
        RECT 101.210 53.770 105.260 54.850 ;
        RECT 66.210 53.020 66.750 53.290 ;
        RECT 67.290 53.020 68.640 53.290 ;
        RECT 69.180 53.020 69.720 53.290 ;
        RECT 83.230 53.030 84.040 53.300 ;
        RECT 84.850 53.030 85.120 53.300 ;
        RECT 85.390 53.030 85.660 53.300 ;
        RECT 85.930 53.030 86.200 53.300 ;
        RECT 86.470 53.030 86.740 53.300 ;
        RECT 87.550 53.030 88.360 53.300 ;
        RECT 101.480 53.230 104.990 53.770 ;
        RECT 66.210 52.750 66.480 53.020 ;
        RECT 65.940 52.480 66.480 52.750 ;
        RECT 65.940 52.210 66.750 52.480 ;
        RECT 67.560 52.210 68.370 53.020 ;
        RECT 69.450 52.750 69.720 53.020 ;
        RECT 69.450 52.480 69.990 52.750 ;
        RECT 84.850 52.490 86.740 53.030 ;
        RECT 102.020 52.960 104.450 53.230 ;
        RECT 105.410 53.210 106.410 53.660 ;
        RECT 106.010 53.110 106.410 53.210 ;
        RECT 102.020 52.690 104.180 52.960 ;
        RECT 69.180 52.210 69.990 52.480 ;
        RECT 65.940 51.130 69.990 52.210 ;
        RECT 84.310 52.220 85.390 52.490 ;
        RECT 86.200 52.220 87.010 52.490 ;
        RECT 84.310 51.950 85.660 52.220 ;
        RECT 85.930 51.950 87.550 52.220 ;
        RECT 84.040 51.680 84.580 51.950 ;
        RECT 85.120 51.680 86.470 51.950 ;
        RECT 87.010 51.680 87.550 51.950 ;
        RECT 84.040 51.410 84.310 51.680 ;
        RECT 83.770 51.140 84.310 51.410 ;
        RECT 66.210 50.590 69.720 51.130 ;
        RECT 66.750 50.320 69.180 50.590 ;
        RECT 70.140 50.570 71.140 51.020 ;
        RECT 70.740 50.470 71.140 50.570 ;
        RECT 83.770 50.870 84.580 51.140 ;
        RECT 85.390 50.870 86.200 51.680 ;
        RECT 87.280 51.410 87.550 51.680 ;
        RECT 87.280 51.140 87.820 51.410 ;
        RECT 87.010 50.870 87.820 51.140 ;
        RECT 66.750 50.050 68.910 50.320 ;
        RECT 83.770 49.790 87.820 50.870 ;
        RECT 84.040 49.250 87.550 49.790 ;
        RECT 84.580 48.980 87.010 49.250 ;
        RECT 87.970 49.230 88.970 49.680 ;
        RECT 88.570 49.130 88.970 49.230 ;
        RECT 84.580 48.710 86.740 48.980 ;
      LAYER met2 ;
        RECT 85.860 223.640 86.180 224.140 ;
        RECT 88.620 223.640 88.940 224.140 ;
        RECT 85.870 222.770 86.130 223.640 ;
        RECT 64.330 222.510 86.130 222.770 ;
        RECT 64.330 219.110 64.590 222.510 ;
        RECT 88.640 222.250 88.900 223.640 ;
        RECT 74.040 221.990 88.900 222.250 ;
        RECT 64.320 218.750 64.630 219.110 ;
        RECT 74.040 219.070 74.300 221.990 ;
        RECT 91.380 221.830 91.700 224.140 ;
        RECT 83.680 221.570 91.700 221.830 ;
        RECT 83.680 219.170 83.940 221.570 ;
        RECT 91.770 220.815 92.250 221.395 ;
        RECT 90.300 219.355 90.760 220.010 ;
        RECT 61.410 218.030 62.100 218.730 ;
        RECT 73.990 218.710 74.300 219.070 ;
        RECT 83.630 218.810 83.940 219.170 ;
        RECT 79.450 187.600 81.440 187.610 ;
        RECT 78.540 187.580 82.340 187.600 ;
        RECT 77.640 187.550 83.240 187.580 ;
        RECT 76.730 187.510 84.150 187.550 ;
        RECT 75.830 187.460 85.050 187.510 ;
        RECT 74.920 187.400 85.960 187.460 ;
        RECT 74.020 187.330 86.860 187.400 ;
        RECT 73.120 187.240 87.760 187.330 ;
        RECT 72.220 187.150 88.660 187.240 ;
        RECT 71.320 187.040 89.560 187.150 ;
        RECT 70.420 186.920 90.460 187.040 ;
        RECT 69.520 186.790 91.360 186.920 ;
        RECT 68.630 186.650 92.250 186.790 ;
        RECT 67.740 186.490 93.140 186.650 ;
        RECT 66.840 186.330 94.040 186.490 ;
        RECT 65.950 186.150 94.930 186.330 ;
        RECT 65.070 185.970 95.810 186.150 ;
        RECT 64.180 185.770 96.700 185.970 ;
        RECT 63.300 185.600 97.580 185.770 ;
        RECT 63.300 185.580 79.640 185.600 ;
        RECT 81.240 185.580 97.580 185.600 ;
        RECT 63.300 185.560 78.730 185.580 ;
        RECT 62.420 185.550 78.730 185.560 ;
        RECT 82.150 185.560 97.580 185.580 ;
        RECT 82.150 185.550 98.460 185.560 ;
        RECT 62.420 185.510 77.830 185.550 ;
        RECT 62.420 185.460 76.920 185.510 ;
        RECT 62.420 185.400 76.020 185.460 ;
        RECT 62.420 185.340 75.120 185.400 ;
        RECT 61.540 185.330 75.120 185.340 ;
        RECT 61.540 185.240 74.220 185.330 ;
        RECT 61.540 185.150 73.320 185.240 ;
        RECT 61.540 185.110 72.420 185.150 ;
        RECT 60.660 185.040 72.420 185.110 ;
        RECT 60.660 184.920 71.520 185.040 ;
        RECT 60.660 184.870 70.630 184.920 ;
        RECT 59.790 184.790 70.630 184.870 ;
        RECT 59.790 184.650 69.740 184.790 ;
        RECT 59.790 184.620 68.840 184.650 ;
        RECT 58.920 184.490 68.840 184.620 ;
        RECT 58.920 184.360 67.950 184.490 ;
        RECT 58.060 184.330 67.950 184.360 ;
        RECT 58.060 184.150 67.070 184.330 ;
        RECT 58.060 184.080 66.180 184.150 ;
        RECT 57.200 183.970 66.180 184.080 ;
        RECT 57.200 183.800 65.300 183.970 ;
        RECT 56.340 183.770 65.300 183.800 ;
        RECT 56.340 183.560 64.420 183.770 ;
        RECT 56.340 183.500 63.540 183.560 ;
        RECT 55.480 183.340 63.540 183.500 ;
        RECT 55.480 183.190 62.660 183.340 ;
        RECT 54.630 183.110 62.660 183.190 ;
        RECT 54.630 182.880 61.790 183.110 ;
        RECT 53.780 182.870 61.790 182.880 ;
        RECT 53.780 182.620 60.920 182.870 ;
        RECT 53.780 182.550 60.060 182.620 ;
        RECT 52.940 182.360 60.060 182.550 ;
        RECT 52.940 182.210 59.200 182.360 ;
        RECT 52.100 182.080 59.200 182.210 ;
        RECT 52.100 181.860 58.340 182.080 ;
        RECT 51.270 181.800 58.340 181.860 ;
        RECT 51.270 181.500 57.480 181.800 ;
        RECT 50.440 181.190 56.630 181.500 ;
        RECT 50.440 181.130 55.780 181.190 ;
        RECT 49.610 180.880 55.780 181.130 ;
        RECT 49.610 180.750 54.940 180.880 ;
        RECT 48.790 180.550 54.940 180.750 ;
        RECT 48.790 180.360 54.100 180.550 ;
        RECT 47.970 180.210 54.100 180.360 ;
        RECT 47.970 179.960 53.270 180.210 ;
        RECT 47.160 179.860 53.270 179.960 ;
        RECT 47.160 179.550 52.440 179.860 ;
        RECT 46.360 179.500 52.440 179.550 ;
        RECT 46.360 179.130 51.610 179.500 ;
        RECT 45.550 178.750 50.790 179.130 ;
        RECT 45.550 178.700 49.970 178.750 ;
        RECT 64.590 178.700 64.990 183.770 ;
        RECT 82.420 180.040 82.820 185.550 ;
        RECT 83.050 185.510 98.460 185.550 ;
        RECT 83.960 185.460 98.460 185.510 ;
        RECT 84.860 185.400 98.460 185.460 ;
        RECT 85.760 185.340 98.460 185.400 ;
        RECT 85.760 185.330 99.340 185.340 ;
        RECT 86.660 185.240 99.340 185.330 ;
        RECT 87.560 185.150 99.340 185.240 ;
        RECT 88.460 185.110 99.340 185.150 ;
        RECT 88.460 185.040 100.220 185.110 ;
        RECT 89.360 184.920 100.220 185.040 ;
        RECT 90.250 184.870 100.220 184.920 ;
        RECT 90.250 184.790 101.090 184.870 ;
        RECT 91.140 184.650 101.090 184.790 ;
        RECT 92.040 184.620 101.090 184.650 ;
        RECT 92.040 184.490 101.960 184.620 ;
        RECT 92.930 184.360 101.960 184.490 ;
        RECT 92.930 184.330 102.820 184.360 ;
        RECT 93.810 184.150 102.820 184.330 ;
        RECT 94.700 184.080 102.820 184.150 ;
        RECT 94.700 183.970 103.680 184.080 ;
        RECT 95.580 183.800 103.680 183.970 ;
        RECT 95.580 183.770 104.540 183.800 ;
        RECT 96.460 183.560 104.540 183.770 ;
        RECT 97.340 183.500 104.540 183.560 ;
        RECT 97.340 183.340 105.400 183.500 ;
        RECT 98.220 183.190 105.400 183.340 ;
        RECT 98.220 183.110 106.250 183.190 ;
        RECT 99.090 182.880 106.250 183.110 ;
        RECT 99.090 182.870 107.100 182.880 ;
        RECT 99.860 182.620 107.100 182.870 ;
        RECT 84.650 180.740 86.810 181.010 ;
        RECT 84.380 180.470 86.810 180.740 ;
        RECT 83.840 179.930 87.350 180.470 ;
        RECT 66.820 179.400 68.980 179.670 ;
        RECT 66.550 179.130 68.980 179.400 ;
        RECT 44.760 178.360 49.970 178.700 ;
        RECT 66.010 178.590 69.520 179.130 ;
        RECT 83.570 178.850 87.620 179.930 ;
        RECT 44.760 178.260 49.160 178.360 ;
        RECT 43.970 177.960 49.160 178.260 ;
        RECT 43.970 177.810 48.360 177.960 ;
        RECT 43.180 177.550 48.360 177.810 ;
        RECT 43.180 177.350 47.550 177.550 ;
        RECT 42.410 177.130 47.550 177.350 ;
        RECT 42.410 176.880 46.760 177.130 ;
        RECT 41.630 176.700 46.760 176.880 ;
        RECT 41.630 176.400 45.970 176.700 ;
        RECT 40.870 176.260 45.970 176.400 ;
        RECT 40.870 175.910 45.180 176.260 ;
        RECT 40.100 175.810 45.180 175.910 ;
        RECT 40.100 175.410 44.410 175.810 ;
        RECT 39.350 175.350 44.410 175.410 ;
        RECT 39.350 174.900 43.630 175.350 ;
        RECT 38.600 174.880 43.630 174.900 ;
        RECT 38.600 174.400 42.870 174.880 ;
        RECT 38.600 174.380 42.100 174.400 ;
        RECT 37.860 173.910 42.100 174.380 ;
        RECT 37.860 173.850 41.350 173.910 ;
        RECT 37.120 173.410 41.350 173.850 ;
        RECT 37.120 173.320 40.600 173.410 ;
        RECT 36.400 172.900 40.600 173.320 ;
        RECT 36.400 172.770 39.860 172.900 ;
        RECT 35.670 172.380 39.860 172.770 ;
        RECT 35.670 172.220 39.120 172.380 ;
        RECT 34.960 171.850 39.120 172.220 ;
        RECT 47.950 172.170 48.350 177.550 ;
        RECT 65.740 177.510 69.790 178.590 ;
        RECT 83.570 178.580 84.380 178.850 ;
        RECT 83.570 178.310 84.110 178.580 ;
        RECT 65.740 177.240 66.550 177.510 ;
        RECT 65.740 176.970 66.280 177.240 ;
        RECT 66.010 176.700 66.280 176.970 ;
        RECT 67.360 176.700 68.170 177.510 ;
        RECT 68.980 177.240 69.790 177.510 ;
        RECT 83.840 178.040 84.110 178.310 ;
        RECT 85.190 178.040 86.000 178.850 ;
        RECT 86.810 178.580 87.620 178.850 ;
        RECT 87.080 178.310 87.620 178.580 ;
        RECT 87.080 178.040 87.350 178.310 ;
        RECT 83.840 177.770 84.380 178.040 ;
        RECT 84.920 177.770 86.270 178.040 ;
        RECT 86.810 177.770 87.350 178.040 ;
        RECT 83.840 177.500 85.460 177.770 ;
        RECT 85.730 177.500 87.080 177.770 ;
        RECT 69.250 176.970 69.790 177.240 ;
        RECT 84.380 177.230 85.190 177.500 ;
        RECT 86.000 177.230 87.080 177.500 ;
        RECT 69.250 176.700 69.520 176.970 ;
        RECT 66.010 176.430 66.550 176.700 ;
        RECT 67.090 176.430 68.440 176.700 ;
        RECT 68.980 176.430 69.520 176.700 ;
        RECT 84.650 176.690 86.540 177.230 ;
        RECT 66.010 176.160 67.630 176.430 ;
        RECT 67.900 176.160 69.250 176.430 ;
        RECT 83.030 176.420 83.840 176.690 ;
        RECT 84.650 176.420 84.920 176.690 ;
        RECT 85.190 176.420 85.460 176.690 ;
        RECT 85.730 176.420 86.000 176.690 ;
        RECT 86.270 176.420 86.540 176.690 ;
        RECT 87.350 176.420 88.160 176.690 ;
        RECT 66.550 175.890 67.360 176.160 ;
        RECT 68.170 175.890 69.250 176.160 ;
        RECT 66.820 175.350 68.710 175.890 ;
        RECT 82.760 175.880 84.110 176.420 ;
        RECT 87.080 175.880 88.430 176.420 ;
        RECT 99.860 176.060 100.260 182.620 ;
        RECT 100.820 182.550 107.100 182.620 ;
        RECT 100.820 182.360 107.940 182.550 ;
        RECT 101.680 182.210 107.940 182.360 ;
        RECT 101.680 182.080 108.780 182.210 ;
        RECT 102.540 181.860 108.780 182.080 ;
        RECT 102.540 181.800 109.610 181.860 ;
        RECT 103.400 181.500 109.610 181.800 ;
        RECT 104.250 181.190 110.440 181.500 ;
        RECT 105.100 181.130 110.440 181.190 ;
        RECT 105.100 180.880 111.270 181.130 ;
        RECT 105.940 180.750 111.270 180.880 ;
        RECT 105.940 180.550 112.090 180.750 ;
        RECT 106.780 180.360 112.090 180.550 ;
        RECT 106.780 180.210 112.910 180.360 ;
        RECT 107.610 179.960 112.910 180.210 ;
        RECT 107.610 179.860 113.720 179.960 ;
        RECT 108.440 179.550 113.720 179.860 ;
        RECT 108.440 179.500 114.520 179.550 ;
        RECT 109.270 179.130 114.520 179.500 ;
        RECT 110.090 178.750 115.330 179.130 ;
        RECT 110.910 178.700 115.330 178.750 ;
        RECT 110.910 178.360 116.120 178.700 ;
        RECT 111.720 178.260 116.120 178.360 ;
        RECT 111.720 177.960 116.910 178.260 ;
        RECT 112.520 177.810 116.910 177.960 ;
        RECT 112.520 177.550 117.700 177.810 ;
        RECT 113.330 177.350 117.700 177.550 ;
        RECT 113.330 177.130 118.470 177.350 ;
        RECT 102.090 176.760 104.250 177.030 ;
        RECT 101.820 176.490 104.250 176.760 ;
        RECT 114.120 176.880 118.470 177.130 ;
        RECT 114.120 176.700 119.250 176.880 ;
        RECT 101.280 175.950 104.790 176.490 ;
        RECT 114.910 176.400 119.250 176.700 ;
        RECT 114.910 176.260 120.010 176.400 ;
        RECT 83.030 175.610 84.650 175.880 ;
        RECT 86.540 175.610 88.160 175.880 ;
        RECT 65.200 175.080 66.010 175.350 ;
        RECT 66.820 175.080 67.090 175.350 ;
        RECT 67.360 175.080 67.630 175.350 ;
        RECT 67.900 175.080 68.170 175.350 ;
        RECT 68.440 175.080 68.710 175.350 ;
        RECT 69.520 175.080 70.330 175.350 ;
        RECT 83.840 175.340 84.920 175.610 ;
        RECT 86.270 175.340 87.350 175.610 ;
        RECT 64.930 174.540 66.280 175.080 ;
        RECT 69.250 174.540 70.600 175.080 ;
        RECT 84.380 175.070 85.460 175.340 ;
        RECT 85.730 175.070 86.810 175.340 ;
        RECT 65.200 174.270 66.820 174.540 ;
        RECT 68.710 174.270 70.330 174.540 ;
        RECT 84.920 174.530 86.270 175.070 ;
        RECT 90.400 174.660 90.740 175.140 ;
        RECT 101.010 174.870 105.060 175.950 ;
        RECT 101.010 174.600 101.820 174.870 ;
        RECT 66.010 174.000 67.090 174.270 ;
        RECT 68.440 174.000 69.520 174.270 ;
        RECT 84.380 174.260 85.460 174.530 ;
        RECT 85.730 174.260 86.810 174.530 ;
        RECT 101.010 174.330 101.550 174.600 ;
        RECT 66.550 173.730 67.630 174.000 ;
        RECT 67.900 173.730 68.980 174.000 ;
        RECT 83.030 173.990 84.920 174.260 ;
        RECT 86.270 173.990 88.430 174.260 ;
        RECT 67.090 173.190 68.440 173.730 ;
        RECT 82.760 173.720 84.380 173.990 ;
        RECT 86.810 173.720 88.430 173.990 ;
        RECT 82.760 173.450 83.840 173.720 ;
        RECT 87.350 173.450 88.430 173.720 ;
        RECT 101.280 174.060 101.550 174.330 ;
        RECT 102.630 174.060 103.440 174.870 ;
        RECT 104.250 174.600 105.060 174.870 ;
        RECT 104.520 174.330 105.060 174.600 ;
        RECT 115.340 175.910 120.010 176.260 ;
        RECT 115.340 175.810 120.780 175.910 ;
        RECT 104.520 174.060 104.790 174.330 ;
        RECT 101.280 173.790 101.820 174.060 ;
        RECT 102.360 173.790 103.710 174.060 ;
        RECT 104.250 173.790 104.790 174.060 ;
        RECT 101.280 173.520 102.900 173.790 ;
        RECT 103.170 173.520 104.520 173.790 ;
        RECT 50.180 172.870 52.340 173.140 ;
        RECT 66.550 172.920 67.630 173.190 ;
        RECT 67.900 172.920 68.980 173.190 ;
        RECT 82.760 173.180 83.570 173.450 ;
        RECT 87.620 173.180 88.430 173.450 ;
        RECT 101.820 173.250 102.630 173.520 ;
        RECT 103.440 173.250 104.520 173.520 ;
        RECT 49.910 172.600 52.340 172.870 ;
        RECT 65.200 172.650 67.090 172.920 ;
        RECT 68.440 172.650 70.600 172.920 ;
        RECT 83.030 172.910 83.300 173.180 ;
        RECT 84.650 172.910 84.920 173.180 ;
        RECT 85.190 172.910 85.460 173.180 ;
        RECT 85.730 172.910 86.000 173.180 ;
        RECT 86.270 172.910 86.540 173.180 ;
        RECT 87.890 172.910 88.160 173.180 ;
        RECT 49.370 172.060 52.880 172.600 ;
        RECT 64.930 172.380 66.550 172.650 ;
        RECT 68.980 172.380 70.600 172.650 ;
        RECT 64.930 172.110 66.010 172.380 ;
        RECT 69.520 172.110 70.600 172.380 ;
        RECT 84.650 172.370 86.540 172.910 ;
        RECT 102.090 172.710 103.980 173.250 ;
        RECT 100.470 172.440 101.280 172.710 ;
        RECT 102.090 172.440 102.360 172.710 ;
        RECT 102.630 172.440 102.900 172.710 ;
        RECT 103.170 172.440 103.440 172.710 ;
        RECT 103.710 172.440 103.980 172.710 ;
        RECT 104.790 172.440 105.600 172.710 ;
        RECT 34.960 171.650 38.400 171.850 ;
        RECT 34.250 171.320 38.400 171.650 ;
        RECT 34.250 171.080 37.670 171.320 ;
        RECT 33.550 170.770 37.670 171.080 ;
        RECT 49.100 170.980 53.150 172.060 ;
        RECT 64.930 171.840 65.740 172.110 ;
        RECT 69.790 171.840 70.600 172.110 ;
        RECT 84.380 172.100 85.190 172.370 ;
        RECT 86.000 172.100 87.080 172.370 ;
        RECT 65.200 171.570 65.470 171.840 ;
        RECT 66.820 171.570 67.090 171.840 ;
        RECT 67.360 171.570 67.630 171.840 ;
        RECT 67.900 171.570 68.170 171.840 ;
        RECT 68.440 171.570 68.710 171.840 ;
        RECT 70.060 171.570 70.330 171.840 ;
        RECT 83.840 171.830 85.460 172.100 ;
        RECT 85.730 171.830 87.080 172.100 ;
        RECT 100.200 171.900 101.550 172.440 ;
        RECT 104.520 171.900 105.870 172.440 ;
        RECT 66.820 171.030 68.710 171.570 ;
        RECT 83.840 171.560 84.380 171.830 ;
        RECT 84.920 171.560 86.270 171.830 ;
        RECT 86.810 171.560 87.350 171.830 ;
        RECT 100.470 171.630 102.090 171.900 ;
        RECT 103.980 171.630 105.600 171.900 ;
        RECT 83.840 171.290 84.110 171.560 ;
        RECT 33.550 170.500 36.960 170.770 ;
        RECT 32.860 170.220 36.960 170.500 ;
        RECT 49.100 170.710 49.910 170.980 ;
        RECT 49.100 170.440 49.640 170.710 ;
        RECT 32.860 169.910 36.250 170.220 ;
        RECT 32.170 169.650 36.250 169.910 ;
        RECT 49.370 170.170 49.640 170.440 ;
        RECT 50.720 170.170 51.530 170.980 ;
        RECT 52.340 170.710 53.150 170.980 ;
        RECT 66.550 170.760 67.360 171.030 ;
        RECT 68.170 170.760 69.250 171.030 ;
        RECT 52.610 170.440 53.150 170.710 ;
        RECT 66.010 170.490 67.630 170.760 ;
        RECT 67.900 170.490 69.250 170.760 ;
        RECT 83.570 171.020 84.110 171.290 ;
        RECT 83.570 170.750 84.380 171.020 ;
        RECT 85.190 170.750 86.000 171.560 ;
        RECT 87.080 171.290 87.350 171.560 ;
        RECT 101.280 171.360 102.360 171.630 ;
        RECT 103.710 171.360 104.790 171.630 ;
        RECT 87.080 171.020 87.620 171.290 ;
        RECT 101.820 171.090 102.900 171.360 ;
        RECT 103.170 171.090 104.250 171.360 ;
        RECT 86.810 170.750 87.620 171.020 ;
        RECT 52.610 170.170 52.880 170.440 ;
        RECT 49.370 169.900 49.910 170.170 ;
        RECT 50.450 169.900 51.800 170.170 ;
        RECT 52.340 169.900 52.880 170.170 ;
        RECT 66.010 170.220 66.550 170.490 ;
        RECT 67.090 170.220 68.440 170.490 ;
        RECT 68.980 170.220 69.520 170.490 ;
        RECT 66.010 169.950 66.280 170.220 ;
        RECT 32.170 169.310 35.550 169.650 ;
        RECT 49.370 169.630 50.990 169.900 ;
        RECT 51.260 169.630 52.610 169.900 ;
        RECT 49.910 169.360 50.720 169.630 ;
        RECT 51.530 169.360 52.610 169.630 ;
        RECT 65.740 169.680 66.280 169.950 ;
        RECT 65.740 169.410 66.550 169.680 ;
        RECT 67.360 169.410 68.170 170.220 ;
        RECT 69.250 169.950 69.520 170.220 ;
        RECT 69.250 169.680 69.790 169.950 ;
        RECT 68.980 169.410 69.790 169.680 ;
        RECT 83.570 169.670 87.620 170.750 ;
        RECT 102.360 170.550 103.710 171.090 ;
        RECT 101.820 170.280 102.900 170.550 ;
        RECT 103.170 170.280 104.250 170.550 ;
        RECT 100.470 170.010 102.360 170.280 ;
        RECT 103.710 170.010 105.870 170.280 ;
        RECT 100.200 169.740 101.820 170.010 ;
        RECT 104.250 169.740 105.870 170.010 ;
        RECT 31.490 169.080 35.550 169.310 ;
        RECT 31.490 168.710 34.860 169.080 ;
        RECT 50.180 168.820 52.070 169.360 ;
        RECT 30.820 168.500 34.860 168.710 ;
        RECT 48.560 168.550 49.370 168.820 ;
        RECT 50.180 168.550 50.450 168.820 ;
        RECT 50.720 168.550 50.990 168.820 ;
        RECT 51.260 168.550 51.530 168.820 ;
        RECT 51.800 168.550 52.070 168.820 ;
        RECT 52.880 168.550 53.690 168.820 ;
        RECT 30.820 168.090 34.360 168.500 ;
        RECT 30.160 167.910 34.360 168.090 ;
        RECT 48.290 168.010 49.640 168.550 ;
        RECT 52.610 168.010 53.960 168.550 ;
        RECT 65.740 168.330 69.790 169.410 ;
        RECT 82.420 168.740 82.920 169.490 ;
        RECT 83.840 169.130 87.350 169.670 ;
        RECT 100.200 169.470 101.280 169.740 ;
        RECT 104.790 169.470 105.870 169.740 ;
        RECT 100.200 169.200 101.010 169.470 ;
        RECT 105.060 169.200 105.870 169.470 ;
        RECT 84.380 168.860 86.810 169.130 ;
        RECT 100.470 168.930 100.740 169.200 ;
        RECT 102.090 168.930 102.360 169.200 ;
        RECT 102.630 168.930 102.900 169.200 ;
        RECT 103.170 168.930 103.440 169.200 ;
        RECT 103.710 168.930 103.980 169.200 ;
        RECT 105.330 168.930 105.600 169.200 ;
        RECT 30.160 167.470 33.490 167.910 ;
        RECT 29.500 167.310 33.490 167.470 ;
        RECT 29.500 166.840 32.820 167.310 ;
        RECT 28.850 166.710 32.820 166.840 ;
        RECT 28.850 166.200 32.160 166.710 ;
        RECT 28.210 166.090 32.160 166.200 ;
        RECT 28.210 165.550 31.500 166.090 ;
        RECT 27.580 165.470 31.500 165.550 ;
        RECT 27.580 164.890 30.850 165.470 ;
        RECT 26.960 164.840 30.850 164.890 ;
        RECT 26.960 164.230 30.210 164.840 ;
        RECT 26.340 164.200 30.210 164.230 ;
        RECT 26.340 163.560 29.580 164.200 ;
        RECT 25.740 163.550 29.580 163.560 ;
        RECT 25.740 162.890 28.960 163.550 ;
        RECT 25.740 162.880 28.340 162.890 ;
        RECT 25.140 162.230 28.340 162.880 ;
        RECT 25.140 162.190 27.740 162.230 ;
        RECT 24.550 161.560 27.740 162.190 ;
        RECT 24.550 161.500 27.140 161.560 ;
        RECT 23.970 160.880 27.140 161.500 ;
        RECT 33.960 161.020 34.360 167.910 ;
        RECT 48.560 167.740 50.180 168.010 ;
        RECT 52.070 167.740 53.690 168.010 ;
        RECT 49.370 167.470 50.450 167.740 ;
        RECT 51.800 167.470 52.880 167.740 ;
        RECT 49.910 167.200 50.990 167.470 ;
        RECT 51.260 167.200 52.340 167.470 ;
        RECT 64.590 167.400 65.090 168.150 ;
        RECT 66.010 167.790 69.520 168.330 ;
        RECT 81.900 168.240 82.920 168.740 ;
        RECT 84.650 168.590 86.810 168.860 ;
        RECT 102.090 168.390 103.980 168.930 ;
        RECT 66.550 167.520 68.980 167.790 ;
        RECT 50.450 166.660 51.800 167.200 ;
        RECT 64.280 166.900 65.090 167.400 ;
        RECT 66.820 167.250 68.980 167.520 ;
        RECT 49.910 166.390 50.990 166.660 ;
        RECT 51.260 166.390 52.340 166.660 ;
        RECT 48.560 166.120 50.450 166.390 ;
        RECT 51.800 166.120 53.960 166.390 ;
        RECT 48.290 165.850 49.910 166.120 ;
        RECT 52.340 165.850 53.960 166.120 ;
        RECT 48.290 165.580 49.370 165.850 ;
        RECT 52.880 165.580 53.960 165.850 ;
        RECT 48.290 165.310 49.100 165.580 ;
        RECT 53.150 165.310 53.960 165.580 ;
        RECT 48.560 165.040 48.830 165.310 ;
        RECT 50.180 165.040 50.450 165.310 ;
        RECT 50.720 165.040 50.990 165.310 ;
        RECT 51.260 165.040 51.530 165.310 ;
        RECT 51.800 165.040 52.070 165.310 ;
        RECT 53.420 165.040 53.690 165.310 ;
        RECT 50.180 164.500 52.070 165.040 ;
        RECT 49.910 164.230 50.720 164.500 ;
        RECT 51.530 164.230 52.610 164.500 ;
        RECT 49.370 163.960 50.990 164.230 ;
        RECT 51.260 163.960 52.610 164.230 ;
        RECT 49.370 163.690 49.910 163.960 ;
        RECT 50.450 163.690 51.800 163.960 ;
        RECT 52.340 163.690 52.880 163.960 ;
        RECT 49.370 163.420 49.640 163.690 ;
        RECT 49.100 163.150 49.640 163.420 ;
        RECT 49.100 162.880 49.910 163.150 ;
        RECT 50.720 162.880 51.530 163.690 ;
        RECT 52.610 163.420 52.880 163.690 ;
        RECT 52.610 163.150 53.150 163.420 ;
        RECT 52.340 162.880 53.150 163.150 ;
        RECT 36.190 161.720 38.350 161.990 ;
        RECT 49.100 161.800 53.150 162.880 ;
        RECT 64.280 162.210 64.780 166.900 ;
        RECT 79.450 164.600 81.440 164.610 ;
        RECT 81.900 164.600 82.400 168.240 ;
        RECT 101.820 168.120 102.630 168.390 ;
        RECT 103.440 168.120 104.520 168.390 ;
        RECT 101.280 167.850 102.900 168.120 ;
        RECT 103.170 167.850 104.520 168.120 ;
        RECT 101.280 167.580 101.820 167.850 ;
        RECT 102.360 167.580 103.710 167.850 ;
        RECT 104.250 167.580 104.790 167.850 ;
        RECT 101.280 167.310 101.550 167.580 ;
        RECT 101.010 167.040 101.550 167.310 ;
        RECT 101.010 166.770 101.820 167.040 ;
        RECT 102.630 166.770 103.440 167.580 ;
        RECT 104.520 167.310 104.790 167.580 ;
        RECT 104.520 167.040 105.060 167.310 ;
        RECT 115.340 167.110 115.740 175.810 ;
        RECT 116.470 175.410 120.780 175.810 ;
        RECT 116.470 175.350 121.530 175.410 ;
        RECT 117.250 174.900 121.530 175.350 ;
        RECT 117.250 174.880 122.280 174.900 ;
        RECT 118.010 174.400 122.280 174.880 ;
        RECT 118.780 174.380 122.280 174.400 ;
        RECT 118.780 173.910 123.020 174.380 ;
        RECT 119.530 173.850 123.020 173.910 ;
        RECT 119.530 173.410 123.760 173.850 ;
        RECT 120.280 173.320 123.760 173.410 ;
        RECT 120.280 172.900 124.480 173.320 ;
        RECT 121.020 172.770 124.480 172.900 ;
        RECT 121.020 172.380 125.210 172.770 ;
        RECT 121.760 172.220 125.210 172.380 ;
        RECT 121.760 171.850 125.920 172.220 ;
        RECT 122.480 171.650 125.920 171.850 ;
        RECT 122.480 171.320 126.630 171.650 ;
        RECT 123.210 171.080 126.630 171.320 ;
        RECT 123.210 170.770 127.330 171.080 ;
        RECT 123.920 170.500 127.330 170.770 ;
        RECT 123.920 170.220 128.020 170.500 ;
        RECT 124.630 169.910 128.020 170.220 ;
        RECT 124.630 169.650 128.710 169.910 ;
        RECT 125.330 169.310 128.710 169.650 ;
        RECT 125.330 169.080 129.390 169.310 ;
        RECT 126.020 168.710 129.390 169.080 ;
        RECT 126.020 168.500 130.060 168.710 ;
        RECT 126.710 168.090 130.060 168.500 ;
        RECT 117.570 167.810 119.730 168.080 ;
        RECT 126.710 167.910 130.720 168.090 ;
        RECT 117.300 167.540 119.730 167.810 ;
        RECT 104.250 166.770 105.060 167.040 ;
        RECT 116.760 167.000 120.270 167.540 ;
        RECT 127.390 167.470 130.720 167.910 ;
        RECT 127.390 167.310 131.380 167.470 ;
        RECT 101.010 165.690 105.060 166.770 ;
        RECT 116.490 165.920 120.540 167.000 ;
        RECT 128.060 166.840 131.380 167.310 ;
        RECT 128.060 166.710 132.030 166.840 ;
        RECT 128.720 166.200 132.030 166.710 ;
        RECT 128.720 166.090 132.670 166.200 ;
        RECT 78.590 164.580 82.400 164.600 ;
        RECT 77.730 164.540 83.150 164.580 ;
        RECT 76.880 164.490 84.000 164.540 ;
        RECT 76.030 164.420 84.850 164.490 ;
        RECT 75.170 164.340 85.710 164.420 ;
        RECT 74.320 164.240 86.560 164.340 ;
        RECT 73.470 164.130 87.410 164.240 ;
        RECT 72.630 164.000 88.250 164.130 ;
        RECT 71.780 163.860 89.100 164.000 ;
        RECT 70.940 163.700 89.940 163.860 ;
        RECT 70.100 163.530 90.780 163.700 ;
        RECT 69.260 163.350 91.620 163.530 ;
        RECT 68.420 163.150 92.460 163.350 ;
        RECT 67.590 162.940 93.290 163.150 ;
        RECT 66.760 162.710 94.120 162.940 ;
        RECT 99.860 162.820 100.360 165.510 ;
        RECT 101.280 165.150 104.790 165.690 ;
        RECT 116.490 165.650 117.300 165.920 ;
        RECT 116.490 165.380 117.030 165.650 ;
        RECT 101.820 164.880 104.250 165.150 ;
        RECT 102.090 164.610 104.250 164.880 ;
        RECT 116.760 165.110 117.030 165.380 ;
        RECT 118.110 165.110 118.920 165.920 ;
        RECT 119.730 165.650 120.540 165.920 ;
        RECT 120.000 165.380 120.540 165.650 ;
        RECT 129.380 165.550 132.670 166.090 ;
        RECT 129.380 165.470 133.300 165.550 ;
        RECT 120.000 165.110 120.270 165.380 ;
        RECT 116.760 164.840 117.300 165.110 ;
        RECT 117.840 164.840 119.190 165.110 ;
        RECT 119.730 164.840 120.270 165.110 ;
        RECT 130.030 164.890 133.300 165.470 ;
        RECT 130.030 164.840 133.920 164.890 ;
        RECT 116.760 164.570 118.380 164.840 ;
        RECT 118.650 164.570 120.000 164.840 ;
        RECT 117.300 164.300 118.110 164.570 ;
        RECT 118.920 164.300 120.000 164.570 ;
        RECT 117.570 163.760 119.460 164.300 ;
        RECT 130.670 164.230 133.920 164.840 ;
        RECT 130.670 164.200 134.540 164.230 ;
        RECT 115.950 163.490 116.760 163.760 ;
        RECT 117.570 163.490 117.840 163.760 ;
        RECT 118.110 163.490 118.380 163.760 ;
        RECT 118.650 163.490 118.920 163.760 ;
        RECT 119.190 163.490 119.460 163.760 ;
        RECT 120.270 163.490 121.080 163.760 ;
        RECT 131.300 163.560 134.540 164.200 ;
        RECT 131.300 163.550 135.140 163.560 ;
        RECT 115.680 162.950 117.030 163.490 ;
        RECT 120.000 162.950 121.350 163.490 ;
        RECT 65.940 162.600 94.940 162.710 ;
        RECT 65.940 162.580 79.730 162.600 ;
        RECT 81.150 162.580 94.940 162.600 ;
        RECT 65.940 162.540 78.880 162.580 ;
        RECT 82.000 162.540 94.940 162.580 ;
        RECT 65.940 162.490 78.030 162.540 ;
        RECT 82.850 162.490 94.940 162.540 ;
        RECT 65.940 162.460 77.170 162.490 ;
        RECT 65.120 162.420 77.170 162.460 ;
        RECT 83.710 162.460 94.940 162.490 ;
        RECT 83.710 162.420 95.760 162.460 ;
        RECT 65.120 162.340 76.320 162.420 ;
        RECT 84.560 162.340 95.760 162.420 ;
        RECT 65.120 162.240 75.470 162.340 ;
        RECT 85.410 162.240 95.760 162.340 ;
        RECT 99.860 162.320 100.700 162.820 ;
        RECT 115.950 162.680 117.570 162.950 ;
        RECT 119.460 162.680 121.080 162.950 ;
        RECT 131.920 162.890 135.140 163.550 ;
        RECT 132.540 162.880 135.140 162.890 ;
        RECT 116.760 162.410 117.840 162.680 ;
        RECT 119.190 162.410 120.270 162.680 ;
        RECT 65.120 162.210 74.630 162.240 ;
        RECT 64.280 162.130 74.630 162.210 ;
        RECT 86.250 162.210 95.760 162.240 ;
        RECT 86.250 162.130 96.580 162.210 ;
        RECT 64.280 162.000 73.780 162.130 ;
        RECT 87.100 162.000 96.580 162.130 ;
        RECT 64.280 161.940 72.940 162.000 ;
        RECT 63.490 161.860 72.940 161.940 ;
        RECT 87.940 161.940 96.580 162.000 ;
        RECT 87.940 161.860 97.390 161.940 ;
        RECT 35.920 161.450 38.350 161.720 ;
        RECT 35.380 160.910 38.890 161.450 ;
        RECT 23.970 160.800 26.550 160.880 ;
        RECT 23.400 160.190 26.550 160.800 ;
        RECT 23.400 160.090 25.970 160.190 ;
        RECT 22.830 159.500 25.970 160.090 ;
        RECT 35.110 159.830 39.160 160.910 ;
        RECT 35.110 159.560 35.920 159.830 ;
        RECT 22.830 159.380 25.400 159.500 ;
        RECT 22.280 158.800 25.400 159.380 ;
        RECT 35.110 159.290 35.650 159.560 ;
        RECT 35.380 159.020 35.650 159.290 ;
        RECT 36.730 159.020 37.540 159.830 ;
        RECT 38.350 159.560 39.160 159.830 ;
        RECT 38.620 159.290 39.160 159.560 ;
        RECT 38.620 159.020 38.890 159.290 ;
        RECT 22.280 158.650 24.830 158.800 ;
        RECT 21.730 158.090 24.830 158.650 ;
        RECT 35.380 158.750 35.920 159.020 ;
        RECT 36.460 158.750 37.810 159.020 ;
        RECT 38.350 158.750 38.890 159.020 ;
        RECT 35.380 158.480 37.000 158.750 ;
        RECT 37.270 158.480 38.620 158.750 ;
        RECT 35.920 158.210 36.730 158.480 ;
        RECT 37.540 158.210 38.620 158.480 ;
        RECT 21.730 157.930 24.280 158.090 ;
        RECT 21.200 157.380 24.280 157.930 ;
        RECT 36.190 157.670 38.080 158.210 ;
        RECT 34.570 157.400 35.380 157.670 ;
        RECT 36.190 157.400 36.460 157.670 ;
        RECT 36.730 157.400 37.000 157.670 ;
        RECT 37.270 157.400 37.540 157.670 ;
        RECT 37.810 157.400 38.080 157.670 ;
        RECT 38.890 157.400 39.700 157.670 ;
        RECT 21.200 157.190 23.730 157.380 ;
        RECT 20.670 156.650 23.730 157.190 ;
        RECT 34.300 156.860 35.650 157.400 ;
        RECT 38.620 156.860 39.970 157.400 ;
        RECT 20.670 156.450 23.200 156.650 ;
        RECT 34.570 156.590 36.190 156.860 ;
        RECT 38.080 156.590 39.700 156.860 ;
        RECT 20.150 155.930 23.200 156.450 ;
        RECT 35.380 156.320 36.460 156.590 ;
        RECT 37.810 156.320 38.890 156.590 ;
        RECT 35.920 156.050 37.000 156.320 ;
        RECT 37.270 156.050 38.350 156.320 ;
        RECT 20.150 155.700 22.670 155.930 ;
        RECT 19.640 155.190 22.670 155.700 ;
        RECT 36.460 155.510 37.810 156.050 ;
        RECT 35.920 155.240 37.000 155.510 ;
        RECT 37.270 155.240 38.350 155.510 ;
        RECT 19.640 154.950 22.150 155.190 ;
        RECT 34.570 154.970 36.460 155.240 ;
        RECT 37.810 154.970 39.970 155.240 ;
        RECT 19.140 154.450 22.150 154.950 ;
        RECT 34.300 154.700 35.920 154.970 ;
        RECT 38.350 154.700 39.970 154.970 ;
        RECT 19.140 154.180 21.640 154.450 ;
        RECT 18.650 153.700 21.640 154.180 ;
        RECT 34.300 154.430 35.380 154.700 ;
        RECT 38.890 154.430 39.970 154.700 ;
        RECT 34.300 154.160 35.110 154.430 ;
        RECT 39.160 154.160 39.970 154.430 ;
        RECT 34.570 153.890 34.840 154.160 ;
        RECT 36.190 153.890 36.460 154.160 ;
        RECT 36.730 153.890 37.000 154.160 ;
        RECT 37.270 153.890 37.540 154.160 ;
        RECT 37.810 153.890 38.080 154.160 ;
        RECT 39.430 153.890 39.700 154.160 ;
        RECT 18.650 153.420 21.140 153.700 ;
        RECT 18.170 152.950 21.140 153.420 ;
        RECT 36.190 153.350 38.080 153.890 ;
        RECT 35.920 153.080 36.730 153.350 ;
        RECT 37.540 153.080 38.620 153.350 ;
        RECT 18.170 152.640 20.650 152.950 ;
        RECT 17.700 152.180 20.650 152.640 ;
        RECT 35.380 152.810 37.000 153.080 ;
        RECT 37.270 152.810 38.620 153.080 ;
        RECT 47.950 153.140 48.450 161.620 ;
        RECT 49.370 161.260 52.880 161.800 ;
        RECT 63.490 161.700 72.100 161.860 ;
        RECT 88.780 161.700 97.390 161.860 ;
        RECT 63.490 161.650 71.260 161.700 ;
        RECT 62.690 161.530 71.260 161.650 ;
        RECT 89.620 161.650 97.390 161.700 ;
        RECT 89.620 161.530 98.190 161.650 ;
        RECT 62.690 161.350 70.420 161.530 ;
        RECT 90.460 161.350 98.190 161.530 ;
        RECT 49.910 160.990 52.340 161.260 ;
        RECT 61.880 161.150 69.590 161.350 ;
        RECT 91.290 161.150 99.000 161.350 ;
        RECT 61.880 161.040 68.760 161.150 ;
        RECT 50.180 160.720 52.340 160.990 ;
        RECT 61.090 160.940 68.760 161.040 ;
        RECT 92.120 161.040 99.000 161.150 ;
        RECT 92.120 160.940 99.790 161.040 ;
        RECT 61.090 160.710 67.940 160.940 ;
        RECT 92.940 160.710 99.790 160.940 ;
        RECT 100.200 160.710 100.700 162.320 ;
        RECT 117.300 162.140 118.380 162.410 ;
        RECT 118.650 162.140 119.730 162.410 ;
        RECT 132.540 162.230 135.740 162.880 ;
        RECT 133.140 162.190 135.740 162.230 ;
        RECT 117.840 161.600 119.190 162.140 ;
        RECT 117.300 161.330 118.380 161.600 ;
        RECT 118.650 161.330 119.730 161.600 ;
        RECT 133.140 161.560 136.330 162.190 ;
        RECT 133.740 161.500 136.330 161.560 ;
        RECT 115.950 161.060 117.840 161.330 ;
        RECT 119.190 161.060 121.350 161.330 ;
        RECT 60.300 160.460 67.120 160.710 ;
        RECT 93.760 160.460 100.700 160.710 ;
        RECT 60.300 160.370 66.300 160.460 ;
        RECT 59.510 160.210 66.300 160.370 ;
        RECT 94.580 160.370 100.700 160.460 ;
        RECT 115.680 160.790 117.300 161.060 ;
        RECT 119.730 160.790 121.350 161.060 ;
        RECT 133.740 160.880 136.910 161.500 ;
        RECT 115.680 160.520 116.760 160.790 ;
        RECT 120.270 160.520 121.350 160.790 ;
        RECT 94.580 160.210 101.370 160.370 ;
        RECT 115.680 160.250 116.490 160.520 ;
        RECT 120.540 160.250 121.350 160.520 ;
        RECT 134.330 160.800 136.910 160.880 ;
        RECT 134.330 160.480 137.480 160.800 ;
        RECT 59.510 160.010 65.490 160.210 ;
        RECT 58.740 159.940 65.490 160.010 ;
        RECT 95.390 160.010 101.370 160.210 ;
        RECT 95.390 159.940 102.140 160.010 ;
        RECT 115.950 159.980 116.220 160.250 ;
        RECT 117.570 159.980 117.840 160.250 ;
        RECT 118.110 159.980 118.380 160.250 ;
        RECT 118.650 159.980 118.920 160.250 ;
        RECT 119.190 159.980 119.460 160.250 ;
        RECT 120.810 159.980 121.080 160.250 ;
        RECT 127.510 160.090 137.480 160.480 ;
        RECT 127.510 160.080 138.050 160.090 ;
        RECT 58.740 159.650 64.690 159.940 ;
        RECT 96.190 159.650 102.140 159.940 ;
        RECT 57.960 159.350 63.880 159.650 ;
        RECT 97.000 159.350 102.920 159.650 ;
        RECT 117.570 159.440 119.460 159.980 ;
        RECT 57.960 159.260 63.090 159.350 ;
        RECT 57.200 159.040 63.090 159.260 ;
        RECT 97.790 159.260 102.920 159.350 ;
        RECT 97.790 159.040 103.680 159.260 ;
        RECT 117.300 159.170 118.110 159.440 ;
        RECT 118.920 159.170 120.000 159.440 ;
        RECT 57.200 158.870 62.300 159.040 ;
        RECT 56.440 158.710 62.300 158.870 ;
        RECT 98.580 158.870 103.680 159.040 ;
        RECT 116.760 158.900 118.380 159.170 ;
        RECT 118.650 158.900 120.000 159.170 ;
        RECT 98.580 158.710 104.440 158.870 ;
        RECT 56.440 158.460 61.510 158.710 ;
        RECT 55.690 158.370 61.510 158.460 ;
        RECT 99.370 158.460 104.440 158.710 ;
        RECT 116.760 158.630 117.300 158.900 ;
        RECT 117.840 158.630 119.190 158.900 ;
        RECT 119.730 158.630 120.270 158.900 ;
        RECT 99.370 158.370 105.190 158.460 ;
        RECT 55.690 158.040 60.740 158.370 ;
        RECT 54.950 158.010 60.740 158.040 ;
        RECT 100.140 158.040 105.190 158.370 ;
        RECT 116.760 158.360 117.030 158.630 ;
        RECT 116.490 158.090 117.030 158.360 ;
        RECT 100.140 158.010 105.940 158.040 ;
        RECT 54.950 157.650 59.960 158.010 ;
        RECT 100.920 157.650 105.940 158.010 ;
        RECT 54.950 157.610 59.200 157.650 ;
        RECT 54.210 157.260 59.200 157.610 ;
        RECT 101.680 157.610 105.940 157.650 ;
        RECT 116.490 157.820 117.300 158.090 ;
        RECT 118.110 157.820 118.920 158.630 ;
        RECT 120.000 158.360 120.270 158.630 ;
        RECT 120.000 158.090 120.540 158.360 ;
        RECT 119.730 157.820 120.540 158.090 ;
        RECT 101.680 157.260 106.670 157.610 ;
        RECT 54.210 157.160 58.440 157.260 ;
        RECT 53.480 156.870 58.440 157.160 ;
        RECT 102.440 157.160 106.670 157.260 ;
        RECT 102.440 156.870 107.400 157.160 ;
        RECT 53.480 156.700 57.690 156.870 ;
        RECT 52.760 156.460 57.690 156.700 ;
        RECT 103.190 156.700 107.400 156.870 ;
        RECT 116.490 156.740 120.540 157.820 ;
        RECT 103.190 156.460 108.120 156.700 ;
        RECT 52.760 156.230 56.950 156.460 ;
        RECT 52.040 156.040 56.950 156.230 ;
        RECT 103.940 156.230 108.120 156.460 ;
        RECT 103.940 156.040 108.840 156.230 ;
        RECT 52.040 155.740 56.210 156.040 ;
        RECT 51.340 155.610 56.210 155.740 ;
        RECT 104.670 155.740 108.840 156.040 ;
        RECT 104.670 155.610 109.540 155.740 ;
        RECT 51.340 155.250 55.480 155.610 ;
        RECT 50.640 155.160 55.480 155.250 ;
        RECT 105.400 155.250 109.540 155.610 ;
        RECT 105.400 155.160 110.240 155.250 ;
        RECT 50.640 154.740 54.760 155.160 ;
        RECT 49.960 154.700 54.760 154.740 ;
        RECT 49.960 154.230 54.040 154.700 ;
        RECT 49.960 154.220 53.340 154.230 ;
        RECT 49.280 153.740 53.340 154.220 ;
        RECT 49.280 153.690 52.640 153.740 ;
        RECT 48.610 153.250 52.640 153.690 ;
        RECT 48.610 153.140 51.960 153.250 ;
        RECT 35.380 152.540 35.920 152.810 ;
        RECT 36.460 152.540 37.810 152.810 ;
        RECT 38.350 152.540 38.890 152.810 ;
        RECT 47.950 152.740 51.960 153.140 ;
        RECT 47.950 152.590 51.280 152.740 ;
        RECT 35.380 152.270 35.650 152.540 ;
        RECT 17.700 151.870 20.170 152.180 ;
        RECT 17.240 151.420 20.170 151.870 ;
        RECT 35.110 152.000 35.650 152.270 ;
        RECT 35.110 151.730 35.920 152.000 ;
        RECT 36.730 151.730 37.540 152.540 ;
        RECT 38.620 152.270 38.890 152.540 ;
        RECT 38.620 152.000 39.160 152.270 ;
        RECT 47.300 152.220 51.280 152.590 ;
        RECT 47.300 152.020 50.610 152.220 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 106.120 154.740 110.240 155.160 ;
        RECT 106.120 154.700 110.920 154.740 ;
        RECT 106.840 154.230 110.920 154.700 ;
        RECT 107.540 154.220 110.920 154.230 ;
        RECT 107.540 153.740 111.600 154.220 ;
        RECT 108.240 153.690 111.600 153.740 ;
        RECT 108.240 153.250 112.270 153.690 ;
        RECT 108.920 153.140 112.270 153.250 ;
        RECT 108.920 152.740 112.930 153.140 ;
        RECT 109.600 152.590 112.930 152.740 ;
        RECT 109.600 152.220 113.580 152.590 ;
        RECT 38.350 151.730 39.160 152.000 ;
        RECT 17.240 151.080 19.700 151.420 ;
        RECT 16.790 150.640 19.700 151.080 ;
        RECT 35.110 150.650 39.160 151.730 ;
        RECT 46.660 151.690 50.610 152.020 ;
        RECT 46.660 151.440 49.950 151.690 ;
        RECT 46.030 151.140 49.950 151.440 ;
        RECT 46.030 150.850 49.300 151.140 ;
        RECT 16.790 150.290 19.240 150.640 ;
        RECT 16.350 149.870 19.240 150.290 ;
        RECT 16.350 149.500 18.790 149.870 ;
        RECT 15.920 149.080 18.790 149.500 ;
        RECT 15.920 148.690 18.350 149.080 ;
        RECT 15.500 148.290 18.350 148.690 ;
        RECT 15.500 147.890 17.920 148.290 ;
        RECT 15.090 147.540 17.920 147.890 ;
        RECT 15.090 147.140 24.290 147.540 ;
        RECT 15.090 147.080 17.500 147.140 ;
        RECT 14.690 146.690 17.500 147.080 ;
        RECT 14.690 146.260 17.090 146.690 ;
        RECT 14.300 145.890 17.090 146.260 ;
        RECT 23.890 146.240 24.290 147.140 ;
        RECT 26.120 146.940 28.280 147.210 ;
        RECT 25.850 146.670 28.280 146.940 ;
        RECT 25.310 146.130 28.820 146.670 ;
        RECT 14.300 145.440 16.690 145.890 ;
        RECT 13.920 145.080 16.690 145.440 ;
        RECT 13.920 144.610 16.300 145.080 ;
        RECT 13.550 144.260 16.300 144.610 ;
        RECT 25.040 145.050 29.090 146.130 ;
        RECT 25.040 144.780 25.850 145.050 ;
        RECT 25.040 144.510 25.580 144.780 ;
        RECT 13.550 143.780 15.920 144.260 ;
        RECT 13.190 143.440 15.920 143.780 ;
        RECT 25.310 144.240 25.580 144.510 ;
        RECT 26.660 144.240 27.470 145.050 ;
        RECT 28.280 144.780 29.090 145.050 ;
        RECT 28.550 144.510 29.090 144.780 ;
        RECT 33.960 145.250 34.460 150.470 ;
        RECT 35.380 150.110 38.890 150.650 ;
        RECT 45.410 150.590 49.300 150.850 ;
        RECT 45.410 150.250 48.660 150.590 ;
        RECT 35.920 149.840 38.350 150.110 ;
        RECT 36.190 149.570 38.350 149.840 ;
        RECT 44.800 150.020 48.660 150.250 ;
        RECT 44.800 149.640 48.030 150.020 ;
        RECT 44.200 149.440 48.030 149.640 ;
        RECT 68.170 149.600 91.570 152.200 ;
        RECT 110.270 152.020 113.580 152.220 ;
        RECT 110.270 151.690 114.220 152.020 ;
        RECT 110.930 151.440 114.220 151.690 ;
        RECT 110.930 151.140 114.850 151.440 ;
        RECT 111.580 150.850 114.850 151.140 ;
        RECT 115.340 150.850 115.840 156.560 ;
        RECT 116.760 156.200 120.270 156.740 ;
        RECT 117.300 155.930 119.730 156.200 ;
        RECT 117.570 155.660 119.730 155.930 ;
        RECT 127.510 154.000 127.910 160.080 ;
        RECT 134.910 159.500 138.050 160.080 ;
        RECT 135.480 159.380 138.050 159.500 ;
        RECT 135.480 158.800 138.600 159.380 ;
        RECT 136.050 158.650 138.600 158.800 ;
        RECT 136.050 158.090 139.150 158.650 ;
        RECT 136.600 157.930 139.150 158.090 ;
        RECT 136.600 157.380 139.680 157.930 ;
        RECT 137.150 157.190 139.680 157.380 ;
        RECT 137.150 156.650 140.210 157.190 ;
        RECT 137.680 156.450 140.210 156.650 ;
        RECT 137.680 155.930 140.730 156.450 ;
        RECT 138.210 155.700 140.730 155.930 ;
        RECT 138.210 155.190 141.240 155.700 ;
        RECT 129.740 154.700 131.900 154.970 ;
        RECT 129.470 154.430 131.900 154.700 ;
        RECT 138.730 154.950 141.240 155.190 ;
        RECT 138.730 154.450 141.740 154.950 ;
        RECT 128.930 153.890 132.440 154.430 ;
        RECT 139.240 154.180 141.740 154.450 ;
        RECT 128.660 152.810 132.710 153.890 ;
        RECT 139.240 153.700 142.230 154.180 ;
        RECT 139.740 153.420 142.230 153.700 ;
        RECT 139.740 152.950 142.710 153.420 ;
        RECT 128.660 152.540 129.470 152.810 ;
        RECT 128.660 152.270 129.200 152.540 ;
        RECT 128.930 152.000 129.200 152.270 ;
        RECT 130.280 152.000 131.090 152.810 ;
        RECT 131.900 152.540 132.710 152.810 ;
        RECT 132.170 152.270 132.710 152.540 ;
        RECT 140.230 152.640 142.710 152.950 ;
        RECT 132.170 152.000 132.440 152.270 ;
        RECT 140.230 152.180 143.180 152.640 ;
        RECT 128.930 151.730 129.470 152.000 ;
        RECT 130.010 151.730 131.360 152.000 ;
        RECT 131.900 151.730 132.440 152.000 ;
        RECT 140.710 151.870 143.180 152.180 ;
        RECT 128.930 151.460 130.550 151.730 ;
        RECT 130.820 151.460 132.170 151.730 ;
        RECT 129.470 151.190 130.280 151.460 ;
        RECT 131.090 151.190 132.170 151.460 ;
        RECT 140.710 151.420 143.640 151.870 ;
        RECT 111.580 150.590 115.840 150.850 ;
        RECT 129.740 150.650 131.630 151.190 ;
        RECT 141.180 151.080 143.640 151.420 ;
        RECT 112.220 150.250 115.840 150.590 ;
        RECT 128.120 150.380 128.930 150.650 ;
        RECT 129.740 150.380 130.010 150.650 ;
        RECT 130.280 150.380 130.550 150.650 ;
        RECT 130.820 150.380 131.090 150.650 ;
        RECT 131.360 150.380 131.630 150.650 ;
        RECT 132.440 150.380 133.250 150.650 ;
        RECT 141.180 150.640 144.090 151.080 ;
        RECT 112.220 150.020 116.080 150.250 ;
        RECT 112.850 149.640 116.080 150.020 ;
        RECT 127.850 149.840 129.200 150.380 ;
        RECT 132.170 149.840 133.520 150.380 ;
        RECT 141.640 150.290 144.090 150.640 ;
        RECT 141.640 149.870 144.530 150.290 ;
        RECT 44.200 149.020 47.410 149.440 ;
        RECT 43.610 148.850 47.410 149.020 ;
        RECT 43.610 148.390 46.800 148.850 ;
        RECT 43.030 148.250 46.800 148.390 ;
        RECT 43.030 147.750 46.200 148.250 ;
        RECT 42.460 147.640 46.200 147.750 ;
        RECT 42.460 147.100 45.610 147.640 ;
        RECT 41.910 147.020 45.610 147.100 ;
        RECT 41.910 146.440 45.030 147.020 ;
        RECT 41.360 146.390 45.030 146.440 ;
        RECT 41.360 145.770 44.460 146.390 ;
        RECT 40.830 145.750 44.460 145.770 ;
        RECT 40.830 145.250 43.910 145.750 ;
        RECT 33.960 145.100 43.910 145.250 ;
        RECT 33.960 144.750 43.360 145.100 ;
        RECT 28.550 144.240 28.820 144.510 ;
        RECT 40.310 144.440 43.360 144.750 ;
        RECT 40.310 144.410 42.830 144.440 ;
        RECT 25.310 143.970 25.850 144.240 ;
        RECT 26.390 143.970 27.740 144.240 ;
        RECT 28.280 143.970 28.820 144.240 ;
        RECT 25.310 143.700 26.930 143.970 ;
        RECT 27.200 143.700 28.550 143.970 ;
        RECT 39.800 143.770 42.830 144.410 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 112.850 149.440 116.680 149.640 ;
        RECT 128.120 149.570 129.740 149.840 ;
        RECT 131.630 149.570 133.250 149.840 ;
        RECT 113.470 149.020 116.680 149.440 ;
        RECT 128.930 149.300 130.010 149.570 ;
        RECT 131.360 149.300 132.440 149.570 ;
        RECT 142.090 149.500 144.530 149.870 ;
        RECT 129.470 149.030 130.550 149.300 ;
        RECT 130.820 149.030 131.900 149.300 ;
        RECT 142.090 149.080 144.960 149.500 ;
        RECT 113.470 148.850 117.270 149.020 ;
        RECT 114.080 148.390 117.270 148.850 ;
        RECT 130.010 148.490 131.360 149.030 ;
        RECT 142.530 148.690 144.960 149.080 ;
        RECT 114.080 148.250 117.850 148.390 ;
        RECT 114.680 147.750 117.850 148.250 ;
        RECT 129.470 148.220 130.550 148.490 ;
        RECT 130.820 148.220 131.900 148.490 ;
        RECT 142.530 148.290 145.380 148.690 ;
        RECT 128.120 147.950 130.010 148.220 ;
        RECT 131.360 147.950 133.520 148.220 ;
        RECT 114.680 147.640 118.420 147.750 ;
        RECT 115.270 147.100 118.420 147.640 ;
        RECT 127.850 147.680 129.470 147.950 ;
        RECT 131.900 147.680 133.520 147.950 ;
        RECT 127.850 147.410 128.930 147.680 ;
        RECT 132.440 147.410 133.520 147.680 ;
        RECT 142.960 147.890 145.380 148.290 ;
        RECT 142.960 147.500 145.790 147.890 ;
        RECT 127.850 147.140 128.660 147.410 ;
        RECT 132.710 147.140 133.520 147.410 ;
        RECT 115.270 147.020 118.970 147.100 ;
        RECT 115.850 146.440 118.970 147.020 ;
        RECT 128.120 146.870 128.390 147.140 ;
        RECT 129.740 146.870 130.010 147.140 ;
        RECT 130.280 146.870 130.550 147.140 ;
        RECT 130.820 146.870 131.090 147.140 ;
        RECT 131.360 146.870 131.630 147.140 ;
        RECT 132.980 146.870 133.250 147.140 ;
        RECT 143.380 147.080 145.790 147.500 ;
        RECT 115.850 146.390 119.520 146.440 ;
        RECT 116.420 145.770 119.520 146.390 ;
        RECT 129.740 146.330 131.630 146.870 ;
        RECT 143.380 146.690 146.190 147.080 ;
        RECT 129.470 146.060 130.280 146.330 ;
        RECT 131.090 146.060 132.170 146.330 ;
        RECT 128.930 145.790 130.550 146.060 ;
        RECT 130.820 145.790 132.170 146.060 ;
        RECT 143.790 146.260 146.190 146.690 ;
        RECT 143.790 145.890 146.580 146.260 ;
        RECT 116.420 145.750 120.050 145.770 ;
        RECT 116.970 145.100 120.050 145.750 ;
        RECT 128.930 145.520 129.470 145.790 ;
        RECT 130.010 145.520 131.360 145.790 ;
        RECT 131.900 145.520 132.440 145.790 ;
        RECT 128.930 145.250 129.200 145.520 ;
        RECT 117.520 145.090 120.050 145.100 ;
        RECT 117.520 144.440 120.570 145.090 ;
        RECT 118.050 144.410 120.570 144.440 ;
        RECT 128.660 144.980 129.200 145.250 ;
        RECT 128.660 144.710 129.470 144.980 ;
        RECT 130.280 144.710 131.090 145.520 ;
        RECT 132.170 145.250 132.440 145.520 ;
        RECT 144.190 145.440 146.580 145.890 ;
        RECT 132.170 144.980 132.710 145.250 ;
        RECT 144.190 145.080 146.960 145.440 ;
        RECT 131.900 144.710 132.710 144.980 ;
        RECT 39.800 143.710 42.310 143.770 ;
        RECT 13.190 142.950 15.550 143.440 ;
        RECT 25.850 143.430 26.660 143.700 ;
        RECT 27.470 143.430 28.550 143.700 ;
        RECT 12.840 142.610 15.550 142.950 ;
        RECT 26.120 142.890 28.010 143.430 ;
        RECT 39.310 143.090 42.310 143.710 ;
        RECT 39.310 143.010 41.800 143.090 ;
        RECT 24.500 142.620 25.310 142.890 ;
        RECT 26.120 142.620 26.390 142.890 ;
        RECT 26.660 142.620 26.930 142.890 ;
        RECT 27.200 142.620 27.470 142.890 ;
        RECT 27.740 142.620 28.010 142.890 ;
        RECT 28.820 142.620 29.630 142.890 ;
        RECT 12.840 142.110 15.190 142.610 ;
        RECT 12.500 141.780 15.190 142.110 ;
        RECT 24.230 142.080 25.580 142.620 ;
        RECT 28.550 142.080 29.900 142.620 ;
        RECT 38.820 142.410 41.800 143.010 ;
        RECT 38.820 142.290 41.310 142.410 ;
        RECT 24.500 141.810 26.120 142.080 ;
        RECT 28.010 141.810 29.630 142.080 ;
        RECT 12.500 141.270 14.840 141.780 ;
        RECT 25.310 141.540 26.390 141.810 ;
        RECT 27.740 141.540 28.820 141.810 ;
        RECT 38.350 141.710 41.310 142.290 ;
        RECT 38.350 141.570 40.820 141.710 ;
        RECT 25.850 141.270 26.930 141.540 ;
        RECT 27.200 141.270 28.280 141.540 ;
        RECT 12.170 140.950 14.840 141.270 ;
        RECT 12.170 140.420 14.500 140.950 ;
        RECT 26.390 140.730 27.740 141.270 ;
        RECT 37.890 141.010 40.820 141.570 ;
        RECT 37.890 140.840 40.350 141.010 ;
        RECT 25.850 140.460 26.930 140.730 ;
        RECT 27.200 140.460 28.280 140.730 ;
        RECT 11.860 140.110 14.500 140.420 ;
        RECT 24.500 140.190 26.390 140.460 ;
        RECT 27.740 140.190 29.900 140.460 ;
        RECT 11.860 139.570 14.170 140.110 ;
        RECT 11.550 139.270 14.170 139.570 ;
        RECT 24.230 139.920 25.850 140.190 ;
        RECT 28.280 139.920 29.900 140.190 ;
        RECT 37.440 140.290 40.350 140.840 ;
        RECT 37.440 140.100 39.890 140.290 ;
        RECT 24.230 139.650 25.310 139.920 ;
        RECT 28.820 139.650 29.900 139.920 ;
        RECT 24.230 139.380 25.040 139.650 ;
        RECT 29.090 139.380 29.900 139.650 ;
        RECT 37.010 139.570 39.890 140.100 ;
        RECT 11.550 138.710 13.860 139.270 ;
        RECT 24.500 139.110 24.770 139.380 ;
        RECT 26.120 139.110 26.390 139.380 ;
        RECT 26.660 139.110 26.930 139.380 ;
        RECT 27.200 139.110 27.470 139.380 ;
        RECT 27.740 139.110 28.010 139.380 ;
        RECT 29.360 139.110 29.630 139.380 ;
        RECT 37.010 139.360 39.440 139.570 ;
        RECT 11.250 138.420 13.860 138.710 ;
        RECT 26.120 138.570 28.010 139.110 ;
        RECT 36.590 138.840 39.440 139.360 ;
        RECT 36.590 138.610 39.010 138.840 ;
        RECT 11.250 137.850 13.550 138.420 ;
        RECT 25.850 138.300 26.660 138.570 ;
        RECT 27.470 138.300 28.550 138.570 ;
        RECT 10.970 137.570 13.550 137.850 ;
        RECT 25.310 138.030 26.930 138.300 ;
        RECT 27.200 138.030 28.550 138.300 ;
        RECT 36.180 138.100 39.010 138.610 ;
        RECT 25.310 137.760 25.850 138.030 ;
        RECT 26.390 137.760 27.740 138.030 ;
        RECT 28.280 137.760 28.820 138.030 ;
        RECT 36.180 137.850 38.590 138.100 ;
        RECT 10.970 136.990 13.250 137.570 ;
        RECT 25.310 137.490 25.580 137.760 ;
        RECT 10.690 136.710 13.250 136.990 ;
        RECT 25.040 137.220 25.580 137.490 ;
        RECT 25.040 136.950 25.850 137.220 ;
        RECT 26.660 136.950 27.470 137.760 ;
        RECT 28.550 137.490 28.820 137.760 ;
        RECT 28.550 137.220 29.090 137.490 ;
        RECT 28.280 136.950 29.090 137.220 ;
        RECT 35.790 137.360 38.590 137.850 ;
        RECT 35.790 137.090 38.180 137.360 ;
        RECT 10.690 136.130 12.970 136.710 ;
        RECT 10.430 135.850 12.970 136.130 ;
        RECT 25.040 135.870 29.090 136.950 ;
        RECT 35.400 136.610 38.180 137.090 ;
        RECT 35.400 136.310 37.790 136.610 ;
        RECT 10.430 135.260 12.690 135.850 ;
        RECT 10.180 134.990 12.690 135.260 ;
        RECT 10.180 134.390 12.430 134.990 ;
        RECT 9.940 134.130 12.430 134.390 ;
        RECT 9.940 133.510 12.180 134.130 ;
        RECT 9.710 133.260 12.180 133.510 ;
        RECT 23.890 133.900 24.390 135.690 ;
        RECT 25.310 135.330 28.820 135.870 ;
        RECT 35.040 135.850 37.790 136.310 ;
        RECT 35.040 135.540 37.400 135.850 ;
        RECT 25.850 135.060 28.280 135.330 ;
        RECT 26.120 134.790 28.280 135.060 ;
        RECT 34.680 135.090 37.400 135.540 ;
        RECT 34.680 134.750 37.040 135.090 ;
        RECT 34.340 134.310 37.040 134.750 ;
        RECT 34.340 133.960 36.680 134.310 ;
        RECT 34.010 133.900 36.680 133.960 ;
        RECT 23.890 133.540 36.680 133.900 ;
        RECT 60.370 134.000 99.370 144.400 ;
        RECT 118.050 143.770 121.080 144.410 ;
        RECT 118.570 143.710 121.080 143.770 ;
        RECT 118.570 143.090 121.570 143.710 ;
        RECT 128.660 143.630 132.710 144.710 ;
        RECT 144.580 144.610 146.960 145.080 ;
        RECT 144.580 144.260 147.330 144.610 ;
        RECT 144.960 143.780 147.330 144.260 ;
        RECT 119.080 143.010 121.570 143.090 ;
        RECT 119.080 142.700 122.060 143.010 ;
        RECT 127.510 142.700 128.010 143.450 ;
        RECT 128.930 143.090 132.440 143.630 ;
        RECT 144.960 143.440 147.690 143.780 ;
        RECT 129.470 142.820 131.900 143.090 ;
        RECT 119.080 142.410 128.010 142.700 ;
        RECT 129.740 142.550 131.900 142.820 ;
        RECT 145.330 142.950 147.690 143.440 ;
        RECT 145.330 142.610 148.040 142.950 ;
        RECT 119.570 142.200 128.010 142.410 ;
        RECT 119.570 141.710 122.530 142.200 ;
        RECT 145.690 142.110 148.040 142.610 ;
        RECT 145.690 141.780 148.380 142.110 ;
        RECT 120.060 141.570 122.530 141.710 ;
        RECT 120.060 141.010 122.990 141.570 ;
        RECT 120.530 140.840 122.990 141.010 ;
        RECT 146.040 141.270 148.380 141.780 ;
        RECT 146.040 140.950 148.710 141.270 ;
        RECT 120.530 140.290 123.440 140.840 ;
        RECT 120.990 140.100 123.440 140.290 ;
        RECT 146.380 140.420 148.710 140.950 ;
        RECT 146.380 140.110 149.020 140.420 ;
        RECT 120.990 139.570 123.870 140.100 ;
        RECT 146.710 139.710 149.020 140.110 ;
        RECT 121.440 139.360 123.870 139.570 ;
        RECT 141.420 139.570 149.020 139.710 ;
        RECT 121.440 138.840 124.290 139.360 ;
        RECT 141.420 139.310 149.330 139.570 ;
        RECT 121.870 138.610 124.290 138.840 ;
        RECT 121.870 138.100 124.700 138.610 ;
        RECT 137.430 138.590 139.590 138.860 ;
        RECT 137.430 138.320 139.860 138.590 ;
        RECT 122.290 137.850 124.700 138.100 ;
        RECT 122.290 137.360 125.090 137.850 ;
        RECT 136.890 137.780 140.400 138.320 ;
        RECT 141.420 137.890 141.820 139.310 ;
        RECT 146.710 139.270 149.330 139.310 ;
        RECT 147.020 138.710 149.330 139.270 ;
        RECT 147.020 138.420 149.630 138.710 ;
        RECT 147.330 137.850 149.630 138.420 ;
        RECT 122.700 137.090 125.090 137.360 ;
        RECT 122.700 136.610 125.480 137.090 ;
        RECT 123.090 136.310 125.480 136.610 ;
        RECT 136.620 136.700 140.670 137.780 ;
        RECT 147.330 137.570 149.910 137.850 ;
        RECT 147.630 136.990 149.910 137.570 ;
        RECT 147.630 136.710 150.190 136.990 ;
        RECT 136.620 136.430 137.430 136.700 ;
        RECT 123.090 135.850 125.840 136.310 ;
        RECT 136.620 136.160 137.160 136.430 ;
        RECT 123.480 135.540 125.840 135.850 ;
        RECT 136.890 135.890 137.160 136.160 ;
        RECT 138.240 135.890 139.050 136.700 ;
        RECT 139.860 136.430 140.670 136.700 ;
        RECT 140.130 136.160 140.670 136.430 ;
        RECT 140.130 135.890 140.400 136.160 ;
        RECT 136.890 135.620 137.430 135.890 ;
        RECT 137.970 135.620 139.320 135.890 ;
        RECT 139.860 135.620 140.400 135.890 ;
        RECT 147.910 136.130 150.190 136.710 ;
        RECT 147.910 135.850 150.450 136.130 ;
        RECT 123.480 135.090 126.200 135.540 ;
        RECT 123.840 134.750 126.200 135.090 ;
        RECT 137.160 135.350 138.510 135.620 ;
        RECT 138.780 135.350 140.400 135.620 ;
        RECT 137.160 135.080 138.240 135.350 ;
        RECT 139.050 135.080 139.860 135.350 ;
        RECT 148.190 135.260 150.450 135.850 ;
        RECT 123.840 134.310 126.540 134.750 ;
        RECT 137.700 134.540 139.590 135.080 ;
        RECT 148.190 134.990 150.700 135.260 ;
        RECT 23.890 133.400 36.340 133.540 ;
        RECT 9.710 132.630 11.940 133.260 ;
        RECT 34.010 133.170 36.340 133.400 ;
        RECT 9.490 132.390 11.940 132.630 ;
        RECT 33.700 132.750 36.340 133.170 ;
        RECT 9.490 131.750 11.710 132.390 ;
        RECT 33.700 132.360 36.010 132.750 ;
        RECT 9.280 131.510 11.710 131.750 ;
        RECT 33.400 131.960 36.010 132.360 ;
        RECT 33.400 131.560 35.700 131.960 ;
        RECT 9.280 131.370 11.490 131.510 ;
        RECT 9.280 130.970 25.170 131.370 ;
        RECT 9.280 130.870 11.490 130.970 ;
        RECT 9.080 130.630 11.490 130.870 ;
        RECT 9.080 129.980 11.280 130.630 ;
        RECT 8.900 129.750 11.280 129.980 ;
        RECT 20.780 129.850 22.940 130.120 ;
        RECT 8.900 129.100 11.080 129.750 ;
        RECT 20.780 129.580 23.210 129.850 ;
        RECT 8.720 128.870 11.080 129.100 ;
        RECT 20.240 129.040 23.750 129.580 ;
        RECT 24.770 129.150 25.170 130.970 ;
        RECT 33.110 131.170 35.700 131.560 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 33.110 130.750 35.400 131.170 ;
        RECT 32.840 130.360 35.400 130.750 ;
        RECT 32.840 129.930 35.110 130.360 ;
        RECT 32.590 129.560 35.110 129.930 ;
        RECT 32.590 129.110 34.840 129.560 ;
        RECT 8.720 128.210 10.900 128.870 ;
        RECT 8.560 127.980 10.900 128.210 ;
        RECT 8.560 127.310 10.720 127.980 ;
        RECT 19.970 127.960 24.020 129.040 ;
        RECT 32.340 128.750 34.840 129.110 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 32.340 128.290 34.590 128.750 ;
        RECT 19.970 127.690 20.780 127.960 ;
        RECT 19.970 127.420 20.510 127.690 ;
        RECT 8.400 127.100 10.720 127.310 ;
        RECT 20.240 127.150 20.510 127.420 ;
        RECT 21.590 127.150 22.400 127.960 ;
        RECT 23.210 127.690 24.020 127.960 ;
        RECT 23.480 127.420 24.020 127.690 ;
        RECT 32.110 127.930 34.590 128.290 ;
        RECT 32.110 127.460 34.340 127.930 ;
        RECT 23.480 127.150 23.750 127.420 ;
        RECT 8.400 126.420 10.560 127.100 ;
        RECT 20.240 126.880 20.780 127.150 ;
        RECT 21.320 126.880 22.670 127.150 ;
        RECT 23.210 126.880 23.750 127.150 ;
        RECT 8.260 126.210 10.560 126.420 ;
        RECT 20.510 126.610 21.860 126.880 ;
        RECT 22.130 126.610 23.750 126.880 ;
        RECT 31.900 127.110 34.340 127.460 ;
        RECT 31.900 126.630 34.110 127.110 ;
        RECT 20.510 126.340 21.590 126.610 ;
        RECT 22.400 126.340 23.210 126.610 ;
        RECT 8.260 125.530 10.400 126.210 ;
        RECT 21.050 125.800 22.940 126.340 ;
        RECT 31.700 126.290 34.110 126.630 ;
        RECT 19.430 125.530 20.240 125.800 ;
        RECT 21.050 125.530 21.320 125.800 ;
        RECT 21.590 125.530 21.860 125.800 ;
        RECT 22.130 125.530 22.400 125.800 ;
        RECT 22.670 125.530 22.940 125.800 ;
        RECT 23.750 125.530 24.560 125.800 ;
        RECT 31.700 125.790 33.900 126.290 ;
        RECT 8.130 125.310 10.400 125.530 ;
        RECT 8.130 124.630 10.260 125.310 ;
        RECT 19.160 124.990 20.510 125.530 ;
        RECT 23.480 124.990 24.830 125.530 ;
        RECT 31.520 125.460 33.900 125.790 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 124.200 133.960 126.540 134.310 ;
        RECT 136.080 134.270 136.890 134.540 ;
        RECT 137.700 134.270 137.970 134.540 ;
        RECT 138.240 134.270 138.510 134.540 ;
        RECT 138.780 134.270 139.050 134.540 ;
        RECT 139.320 134.270 139.590 134.540 ;
        RECT 140.400 134.270 141.210 134.540 ;
        RECT 148.450 134.390 150.700 134.990 ;
        RECT 124.200 133.540 126.870 133.960 ;
        RECT 135.810 133.730 137.160 134.270 ;
        RECT 140.130 133.730 141.480 134.270 ;
        RECT 148.450 134.130 150.940 134.390 ;
        RECT 124.540 133.170 126.870 133.540 ;
        RECT 136.080 133.460 137.700 133.730 ;
        RECT 139.590 133.460 141.210 133.730 ;
        RECT 148.700 133.510 150.940 134.130 ;
        RECT 136.890 133.190 137.970 133.460 ;
        RECT 139.320 133.190 140.400 133.460 ;
        RECT 148.700 133.260 151.170 133.510 ;
        RECT 124.540 132.750 127.180 133.170 ;
        RECT 137.430 132.920 138.510 133.190 ;
        RECT 138.780 132.920 139.860 133.190 ;
        RECT 124.870 132.360 127.180 132.750 ;
        RECT 137.970 132.380 139.320 132.920 ;
        RECT 148.940 132.630 151.170 133.260 ;
        RECT 148.940 132.390 151.390 132.630 ;
        RECT 124.870 131.960 127.480 132.360 ;
        RECT 137.430 132.110 138.510 132.380 ;
        RECT 138.780 132.110 139.860 132.380 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 125.180 131.560 127.480 131.960 ;
        RECT 135.810 131.840 137.970 132.110 ;
        RECT 139.320 131.840 141.210 132.110 ;
        RECT 135.810 131.570 137.430 131.840 ;
        RECT 139.860 131.570 141.480 131.840 ;
        RECT 125.180 131.170 127.770 131.560 ;
        RECT 125.480 130.750 127.770 131.170 ;
        RECT 135.810 131.300 136.890 131.570 ;
        RECT 140.400 131.300 141.480 131.570 ;
        RECT 149.170 131.750 151.390 132.390 ;
        RECT 149.170 131.510 151.600 131.750 ;
        RECT 135.810 131.030 136.620 131.300 ;
        RECT 140.670 131.030 141.480 131.300 ;
        RECT 136.080 130.760 136.350 131.030 ;
        RECT 137.700 130.760 137.970 131.030 ;
        RECT 138.240 130.760 138.510 131.030 ;
        RECT 138.780 130.760 139.050 131.030 ;
        RECT 139.320 130.760 139.590 131.030 ;
        RECT 140.940 130.760 141.210 131.030 ;
        RECT 149.390 130.870 151.600 131.510 ;
        RECT 125.480 130.360 128.040 130.750 ;
        RECT 125.770 129.930 128.040 130.360 ;
        RECT 137.700 130.220 139.590 130.760 ;
        RECT 149.390 130.630 151.800 130.870 ;
        RECT 137.160 129.950 138.240 130.220 ;
        RECT 139.050 129.950 139.860 130.220 ;
        RECT 149.600 129.980 151.800 130.630 ;
        RECT 125.770 129.560 128.290 129.930 ;
        RECT 137.160 129.680 138.510 129.950 ;
        RECT 138.780 129.680 140.400 129.950 ;
        RECT 149.600 129.750 151.980 129.980 ;
        RECT 126.040 129.110 128.290 129.560 ;
        RECT 136.890 129.410 137.430 129.680 ;
        RECT 137.970 129.410 139.320 129.680 ;
        RECT 139.860 129.410 140.400 129.680 ;
        RECT 136.890 129.140 137.160 129.410 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 126.040 128.750 128.540 129.110 ;
        RECT 126.290 128.290 128.540 128.750 ;
        RECT 136.620 128.870 137.160 129.140 ;
        RECT 136.620 128.600 137.430 128.870 ;
        RECT 138.240 128.600 139.050 129.410 ;
        RECT 140.130 129.140 140.400 129.410 ;
        RECT 140.130 128.870 140.670 129.140 ;
        RECT 149.800 129.100 151.980 129.750 ;
        RECT 149.800 128.870 152.160 129.100 ;
        RECT 139.860 128.600 140.670 128.870 ;
        RECT 126.290 127.930 128.770 128.290 ;
        RECT 126.540 127.460 128.770 127.930 ;
        RECT 136.620 127.520 140.670 128.600 ;
        RECT 149.980 128.210 152.160 128.870 ;
        RECT 149.980 127.980 152.320 128.210 ;
        RECT 126.540 127.110 128.980 127.460 ;
        RECT 126.770 126.630 128.980 127.110 ;
        RECT 136.890 126.980 140.400 127.520 ;
        RECT 137.430 126.710 139.860 126.980 ;
        RECT 126.770 126.290 129.180 126.630 ;
        RECT 137.430 126.440 139.590 126.710 ;
        RECT 19.430 124.720 21.050 124.990 ;
        RECT 22.940 124.720 24.560 124.990 ;
        RECT 31.520 124.950 33.700 125.460 ;
        RECT 8.010 124.420 10.260 124.630 ;
        RECT 20.240 124.450 21.320 124.720 ;
        RECT 22.670 124.450 23.750 124.720 ;
        RECT 31.350 124.630 33.700 124.950 ;
        RECT 8.010 123.730 10.130 124.420 ;
        RECT 20.780 124.180 21.860 124.450 ;
        RECT 22.130 124.180 23.210 124.450 ;
        RECT 7.900 123.530 10.130 123.730 ;
        RECT 21.320 123.640 22.670 124.180 ;
        RECT 31.350 124.110 33.520 124.630 ;
        RECT 31.190 123.790 33.520 124.110 ;
        RECT 7.900 122.830 10.010 123.530 ;
        RECT 20.780 123.370 21.860 123.640 ;
        RECT 22.130 123.370 23.210 123.640 ;
        RECT 7.810 122.630 10.010 122.830 ;
        RECT 19.160 123.100 21.320 123.370 ;
        RECT 22.670 123.100 24.560 123.370 ;
        RECT 31.190 123.270 33.350 123.790 ;
        RECT 19.160 122.830 20.780 123.100 ;
        RECT 23.210 122.830 24.830 123.100 ;
        RECT 7.810 121.930 9.900 122.630 ;
        RECT 19.160 122.560 20.240 122.830 ;
        RECT 23.750 122.560 24.830 122.830 ;
        RECT 19.160 122.290 19.970 122.560 ;
        RECT 24.020 122.290 24.830 122.560 ;
        RECT 31.050 122.950 33.350 123.270 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
        RECT 126.980 125.790 129.180 126.290 ;
        RECT 126.980 125.460 129.360 125.790 ;
        RECT 127.180 125.450 129.360 125.460 ;
        RECT 141.320 125.450 141.820 127.340 ;
        RECT 150.160 127.310 152.320 127.980 ;
        RECT 150.160 127.100 152.480 127.310 ;
        RECT 150.320 126.420 152.480 127.100 ;
        RECT 150.320 126.210 152.620 126.420 ;
        RECT 127.180 124.950 141.820 125.450 ;
        RECT 150.480 125.530 152.620 126.210 ;
        RECT 150.480 125.310 152.750 125.530 ;
        RECT 127.180 124.630 129.530 124.950 ;
        RECT 127.360 124.110 129.530 124.630 ;
        RECT 150.620 124.630 152.750 125.310 ;
        RECT 150.620 124.420 152.870 124.630 ;
        RECT 127.360 123.790 129.690 124.110 ;
        RECT 31.050 122.420 33.190 122.950 ;
        RECT 19.430 122.020 19.700 122.290 ;
        RECT 21.050 122.020 21.320 122.290 ;
        RECT 21.590 122.020 21.860 122.290 ;
        RECT 22.130 122.020 22.400 122.290 ;
        RECT 22.670 122.020 22.940 122.290 ;
        RECT 24.290 122.020 24.560 122.290 ;
        RECT 30.920 122.110 33.190 122.420 ;
        RECT 7.720 121.730 9.900 121.930 ;
        RECT 7.720 121.030 9.810 121.730 ;
        RECT 21.050 121.480 22.940 122.020 ;
        RECT 30.920 121.580 33.050 122.110 ;
        RECT 7.650 120.830 9.810 121.030 ;
        RECT 20.510 121.210 21.590 121.480 ;
        RECT 22.400 121.210 23.210 121.480 ;
        RECT 30.810 121.270 33.050 121.580 ;
        RECT 20.510 120.940 21.860 121.210 ;
        RECT 22.130 120.940 23.750 121.210 ;
        RECT 7.650 120.130 9.720 120.830 ;
        RECT 20.240 120.670 20.780 120.940 ;
        RECT 21.320 120.670 22.670 120.940 ;
        RECT 23.210 120.670 23.750 120.940 ;
        RECT 30.810 120.730 32.920 121.270 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 127.530 123.270 129.690 123.790 ;
        RECT 150.750 123.730 152.870 124.420 ;
        RECT 150.750 123.530 152.980 123.730 ;
        RECT 127.530 122.950 129.830 123.270 ;
        RECT 127.690 122.420 129.830 122.950 ;
        RECT 150.870 122.830 152.980 123.530 ;
        RECT 150.870 122.630 153.070 122.830 ;
        RECT 127.690 122.110 129.960 122.420 ;
        RECT 150.980 122.390 153.070 122.630 ;
        RECT 127.830 121.580 129.960 122.110 ;
        RECT 137.940 121.990 153.070 122.390 ;
        RECT 127.830 121.270 130.070 121.580 ;
        RECT 20.240 120.400 20.510 120.670 ;
        RECT 7.590 119.930 9.720 120.130 ;
        RECT 19.970 120.130 20.510 120.400 ;
        RECT 7.590 119.220 9.650 119.930 ;
        RECT 7.540 119.030 9.650 119.220 ;
        RECT 19.970 119.860 20.780 120.130 ;
        RECT 21.590 119.860 22.400 120.670 ;
        RECT 23.480 120.400 23.750 120.670 ;
        RECT 30.710 120.420 32.920 120.730 ;
        RECT 23.480 120.130 24.020 120.400 ;
        RECT 23.210 119.860 24.020 120.130 ;
        RECT 30.710 119.880 32.810 120.420 ;
        RECT 7.540 118.320 9.590 119.030 ;
        RECT 19.970 118.780 24.020 119.860 ;
        RECT 30.630 119.580 32.810 119.880 ;
        RECT 30.630 119.020 32.710 119.580 ;
        RECT 7.500 118.130 9.590 118.320 ;
        RECT 20.240 118.240 23.750 118.780 ;
        RECT 30.560 118.730 32.710 119.020 ;
        RECT 7.500 117.410 9.540 118.130 ;
        RECT 20.780 117.970 23.210 118.240 ;
        RECT 20.780 117.700 22.940 117.970 ;
        RECT 7.470 117.220 9.540 117.410 ;
        RECT 24.670 117.520 25.170 118.600 ;
        RECT 30.560 118.170 32.630 118.730 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 127.960 120.730 130.070 121.270 ;
        RECT 127.960 120.420 130.170 120.730 ;
        RECT 128.070 119.880 130.170 120.420 ;
        RECT 137.940 120.210 138.340 121.990 ;
        RECT 150.980 121.930 153.070 121.990 ;
        RECT 150.980 121.730 153.160 121.930 ;
        RECT 140.170 120.910 142.330 121.180 ;
        RECT 139.900 120.640 142.330 120.910 ;
        RECT 151.070 121.030 153.160 121.730 ;
        RECT 151.070 120.830 153.230 121.030 ;
        RECT 139.360 120.100 142.870 120.640 ;
        RECT 151.160 120.130 153.230 120.830 ;
        RECT 128.070 119.580 130.250 119.880 ;
        RECT 128.170 119.020 130.250 119.580 ;
        RECT 139.090 119.020 143.140 120.100 ;
        RECT 151.160 119.930 153.290 120.130 ;
        RECT 151.230 119.220 153.290 119.930 ;
        RECT 151.230 119.030 153.340 119.220 ;
        RECT 128.170 118.730 130.320 119.020 ;
        RECT 30.510 117.880 32.630 118.170 ;
        RECT 30.510 117.520 32.560 117.880 ;
        RECT 7.470 116.510 9.500 117.220 ;
        RECT 24.670 117.020 32.560 117.520 ;
        RECT 7.450 116.320 9.500 116.510 ;
        RECT 30.470 116.460 32.510 117.020 ;
        RECT 7.450 115.610 9.470 116.320 ;
        RECT 30.450 116.170 32.510 116.460 ;
        RECT 30.450 115.610 32.470 116.170 ;
        RECT 7.440 115.410 9.470 115.610 ;
        RECT 7.440 113.810 9.450 115.410 ;
        RECT 30.440 115.320 32.470 115.610 ;
        RECT 30.440 113.900 32.450 115.320 ;
        RECT 7.440 113.620 9.470 113.810 ;
        RECT 30.440 113.620 32.470 113.900 ;
        RECT 7.450 112.900 9.470 113.620 ;
        RECT 30.450 113.050 32.470 113.620 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 128.250 118.170 130.320 118.730 ;
        RECT 139.090 118.750 139.900 119.020 ;
        RECT 139.090 118.480 139.630 118.750 ;
        RECT 139.360 118.210 139.630 118.480 ;
        RECT 140.710 118.210 141.520 119.020 ;
        RECT 142.330 118.750 143.140 119.020 ;
        RECT 142.600 118.480 143.140 118.750 ;
        RECT 142.600 118.210 142.870 118.480 ;
        RECT 128.250 117.880 130.370 118.170 ;
        RECT 128.320 117.320 130.370 117.880 ;
        RECT 139.360 117.940 139.900 118.210 ;
        RECT 140.440 117.940 141.790 118.210 ;
        RECT 142.330 117.940 142.870 118.210 ;
        RECT 151.290 118.320 153.340 119.030 ;
        RECT 151.290 118.130 153.380 118.320 ;
        RECT 139.360 117.670 140.980 117.940 ;
        RECT 141.250 117.670 142.600 117.940 ;
        RECT 139.900 117.400 140.710 117.670 ;
        RECT 141.520 117.400 142.600 117.670 ;
        RECT 151.340 117.410 153.380 118.130 ;
        RECT 128.320 117.020 130.410 117.320 ;
        RECT 128.370 116.460 130.410 117.020 ;
        RECT 140.170 116.860 142.060 117.400 ;
        RECT 151.340 117.220 153.410 117.410 ;
        RECT 138.550 116.590 139.360 116.860 ;
        RECT 140.170 116.590 140.440 116.860 ;
        RECT 140.710 116.590 140.980 116.860 ;
        RECT 141.250 116.590 141.520 116.860 ;
        RECT 141.790 116.590 142.060 116.860 ;
        RECT 142.870 116.590 143.680 116.860 ;
        RECT 128.370 116.170 130.430 116.460 ;
        RECT 128.410 115.610 130.430 116.170 ;
        RECT 138.280 116.050 139.630 116.590 ;
        RECT 142.600 116.050 143.950 116.590 ;
        RECT 151.380 116.510 153.410 117.220 ;
        RECT 151.380 116.320 153.430 116.510 ;
        RECT 138.550 115.780 140.170 116.050 ;
        RECT 142.060 115.780 143.680 116.050 ;
        RECT 128.410 115.320 130.440 115.610 ;
        RECT 139.360 115.510 140.440 115.780 ;
        RECT 141.790 115.510 142.870 115.780 ;
        RECT 151.410 115.610 153.430 116.320 ;
        RECT 128.430 113.900 130.440 115.320 ;
        RECT 139.900 115.240 140.980 115.510 ;
        RECT 141.250 115.240 142.330 115.510 ;
        RECT 151.410 115.410 153.440 115.610 ;
        RECT 140.440 114.700 141.790 115.240 ;
        RECT 139.900 114.430 140.980 114.700 ;
        RECT 141.250 114.430 142.330 114.700 ;
        RECT 138.550 114.160 140.440 114.430 ;
        RECT 141.790 114.160 143.950 114.430 ;
        RECT 128.410 113.610 130.440 113.900 ;
        RECT 138.280 113.890 139.900 114.160 ;
        RECT 142.330 113.890 143.950 114.160 ;
        RECT 138.280 113.620 139.360 113.890 ;
        RECT 142.870 113.620 143.950 113.890 ;
        RECT 151.430 113.810 153.440 115.410 ;
        RECT 7.450 112.710 9.500 112.900 ;
        RECT 30.450 112.760 32.510 113.050 ;
        RECT 7.470 112.570 9.500 112.710 ;
        RECT 7.470 112.170 19.020 112.570 ;
        RECT 7.470 112.000 9.500 112.170 ;
        RECT 7.470 111.810 9.540 112.000 ;
        RECT 7.500 111.090 9.540 111.810 ;
        RECT 18.620 111.270 19.020 112.170 ;
        RECT 20.850 111.970 23.010 112.240 ;
        RECT 20.580 111.700 23.010 111.970 ;
        RECT 30.470 112.200 32.510 112.760 ;
        RECT 30.470 111.900 32.560 112.200 ;
        RECT 20.040 111.160 23.550 111.700 ;
        RECT 30.510 111.340 32.560 111.900 ;
        RECT 7.500 110.900 9.590 111.090 ;
        RECT 7.540 110.190 9.590 110.900 ;
        RECT 7.540 110.000 9.650 110.190 ;
        RECT 7.590 109.290 9.650 110.000 ;
        RECT 19.770 110.080 23.820 111.160 ;
        RECT 30.510 111.050 32.630 111.340 ;
        RECT 30.560 110.490 32.630 111.050 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 128.410 113.050 130.430 113.610 ;
        RECT 138.280 113.350 139.090 113.620 ;
        RECT 143.140 113.350 143.950 113.620 ;
        RECT 151.410 113.610 153.440 113.810 ;
        RECT 138.550 113.080 138.820 113.350 ;
        RECT 140.170 113.080 140.440 113.350 ;
        RECT 140.710 113.080 140.980 113.350 ;
        RECT 141.250 113.080 141.520 113.350 ;
        RECT 141.790 113.080 142.060 113.350 ;
        RECT 143.410 113.080 143.680 113.350 ;
        RECT 128.370 112.760 130.430 113.050 ;
        RECT 128.370 112.200 130.410 112.760 ;
        RECT 140.170 112.540 142.060 113.080 ;
        RECT 151.410 112.900 153.430 113.610 ;
        RECT 151.380 112.710 153.430 112.900 ;
        RECT 139.900 112.270 140.710 112.540 ;
        RECT 141.520 112.270 142.600 112.540 ;
        RECT 128.320 111.900 130.410 112.200 ;
        RECT 139.360 112.000 140.980 112.270 ;
        RECT 141.250 112.000 142.600 112.270 ;
        RECT 151.380 112.000 153.410 112.710 ;
        RECT 128.320 111.340 130.370 111.900 ;
        RECT 139.360 111.730 139.900 112.000 ;
        RECT 140.440 111.730 141.790 112.000 ;
        RECT 142.330 111.730 142.870 112.000 ;
        RECT 139.360 111.460 139.630 111.730 ;
        RECT 128.250 111.050 130.370 111.340 ;
        RECT 139.090 111.190 139.630 111.460 ;
        RECT 30.560 110.200 32.710 110.490 ;
        RECT 19.770 109.810 20.580 110.080 ;
        RECT 19.770 109.540 20.310 109.810 ;
        RECT 7.590 109.090 9.720 109.290 ;
        RECT 7.650 108.390 9.720 109.090 ;
        RECT 20.040 109.270 20.310 109.540 ;
        RECT 21.390 109.270 22.200 110.080 ;
        RECT 23.010 109.810 23.820 110.080 ;
        RECT 23.280 109.540 23.820 109.810 ;
        RECT 30.630 109.640 32.710 110.200 ;
        RECT 23.280 109.270 23.550 109.540 ;
        RECT 30.630 109.340 32.810 109.640 ;
        RECT 20.040 109.000 20.580 109.270 ;
        RECT 21.120 109.000 22.470 109.270 ;
        RECT 23.010 109.000 23.550 109.270 ;
        RECT 20.040 108.730 21.660 109.000 ;
        RECT 21.930 108.730 23.280 109.000 ;
        RECT 20.580 108.460 21.390 108.730 ;
        RECT 22.200 108.460 23.280 108.730 ;
        RECT 30.710 108.800 32.810 109.340 ;
        RECT 30.710 108.490 32.920 108.800 ;
        RECT 7.650 108.190 9.810 108.390 ;
        RECT 7.720 107.490 9.810 108.190 ;
        RECT 20.850 107.920 22.740 108.460 ;
        RECT 30.810 107.950 32.920 108.490 ;
        RECT 19.230 107.650 20.040 107.920 ;
        RECT 20.850 107.650 21.120 107.920 ;
        RECT 21.390 107.650 21.660 107.920 ;
        RECT 21.930 107.650 22.200 107.920 ;
        RECT 22.470 107.650 22.740 107.920 ;
        RECT 23.550 107.650 24.360 107.920 ;
        RECT 7.720 107.290 9.900 107.490 ;
        RECT 7.810 106.590 9.900 107.290 ;
        RECT 18.960 107.110 20.310 107.650 ;
        RECT 23.280 107.110 24.630 107.650 ;
        RECT 30.810 107.640 33.050 107.950 ;
        RECT 30.920 107.110 33.050 107.640 ;
        RECT 19.230 106.840 20.850 107.110 ;
        RECT 22.740 106.840 24.360 107.110 ;
        RECT 7.810 106.390 10.010 106.590 ;
        RECT 20.040 106.570 21.120 106.840 ;
        RECT 22.470 106.570 23.550 106.840 ;
        RECT 30.920 106.800 33.190 107.110 ;
        RECT 7.900 105.690 10.010 106.390 ;
        RECT 20.580 106.300 21.660 106.570 ;
        RECT 21.930 106.300 23.010 106.570 ;
        RECT 21.120 105.760 22.470 106.300 ;
        RECT 31.050 106.270 33.190 106.800 ;
        RECT 31.050 105.950 33.350 106.270 ;
        RECT 7.900 105.490 10.130 105.690 ;
        RECT 20.580 105.490 21.660 105.760 ;
        RECT 21.930 105.490 23.010 105.760 ;
        RECT 8.010 104.800 10.130 105.490 ;
        RECT 19.230 105.220 21.120 105.490 ;
        RECT 22.470 105.220 24.630 105.490 ;
        RECT 18.960 104.950 20.580 105.220 ;
        RECT 23.010 104.950 24.630 105.220 ;
        RECT 31.190 105.430 33.350 105.950 ;
        RECT 31.190 105.110 33.520 105.430 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
        RECT 128.250 110.490 130.320 111.050 ;
        RECT 128.170 110.200 130.320 110.490 ;
        RECT 139.090 110.920 139.900 111.190 ;
        RECT 140.710 110.920 141.520 111.730 ;
        RECT 142.600 111.460 142.870 111.730 ;
        RECT 151.340 111.810 153.410 112.000 ;
        RECT 142.600 111.190 143.140 111.460 ;
        RECT 142.330 110.920 143.140 111.190 ;
        RECT 151.340 111.090 153.380 111.810 ;
        RECT 128.170 109.640 130.250 110.200 ;
        RECT 139.090 109.840 143.140 110.920 ;
        RECT 151.290 110.900 153.380 111.090 ;
        RECT 151.290 110.190 153.340 110.900 ;
        RECT 151.230 110.000 153.340 110.190 ;
        RECT 128.070 109.340 130.250 109.640 ;
        RECT 128.070 108.910 130.170 109.340 ;
        RECT 137.940 108.910 138.440 109.660 ;
        RECT 139.360 109.300 142.870 109.840 ;
        RECT 139.900 109.030 142.330 109.300 ;
        RECT 151.230 109.290 153.290 110.000 ;
        RECT 128.070 108.800 138.440 108.910 ;
        RECT 127.960 108.410 138.440 108.800 ;
        RECT 140.170 108.760 142.330 109.030 ;
        RECT 151.160 109.090 153.290 109.290 ;
        RECT 127.960 107.950 130.070 108.410 ;
        RECT 151.160 108.390 153.230 109.090 ;
        RECT 127.830 107.640 130.070 107.950 ;
        RECT 151.070 108.190 153.230 108.390 ;
        RECT 127.830 107.110 129.960 107.640 ;
        RECT 151.070 107.490 153.160 108.190 ;
        RECT 127.690 106.800 129.960 107.110 ;
        RECT 150.980 107.290 153.160 107.490 ;
        RECT 127.690 106.270 129.830 106.800 ;
        RECT 150.980 106.590 153.070 107.290 ;
        RECT 127.530 105.950 129.830 106.270 ;
        RECT 150.870 106.390 153.070 106.590 ;
        RECT 127.530 105.430 129.690 105.950 ;
        RECT 150.870 105.690 152.980 106.390 ;
        RECT 8.010 104.590 10.260 104.800 ;
        RECT 8.130 103.910 10.260 104.590 ;
        RECT 18.960 104.680 20.040 104.950 ;
        RECT 23.550 104.680 24.630 104.950 ;
        RECT 18.960 104.410 19.770 104.680 ;
        RECT 23.820 104.410 24.630 104.680 ;
        RECT 31.350 104.590 33.520 105.110 ;
        RECT 19.230 104.140 19.500 104.410 ;
        RECT 20.850 104.140 21.120 104.410 ;
        RECT 21.390 104.140 21.660 104.410 ;
        RECT 21.930 104.140 22.200 104.410 ;
        RECT 22.470 104.140 22.740 104.410 ;
        RECT 24.090 104.140 24.360 104.410 ;
        RECT 31.350 104.270 33.700 104.590 ;
        RECT 8.130 103.690 10.400 103.910 ;
        RECT 8.260 103.010 10.400 103.690 ;
        RECT 20.850 103.600 22.740 104.140 ;
        RECT 31.520 103.760 33.700 104.270 ;
        RECT 20.580 103.330 21.390 103.600 ;
        RECT 22.200 103.330 23.280 103.600 ;
        RECT 31.520 103.430 33.900 103.760 ;
        RECT 20.040 103.060 21.660 103.330 ;
        RECT 21.930 103.060 23.280 103.330 ;
        RECT 8.260 102.800 10.560 103.010 ;
        RECT 8.400 102.120 10.560 102.800 ;
        RECT 20.040 102.790 20.580 103.060 ;
        RECT 21.120 102.790 22.470 103.060 ;
        RECT 23.010 102.790 23.550 103.060 ;
        RECT 20.040 102.520 20.310 102.790 ;
        RECT 19.770 102.250 20.310 102.520 ;
        RECT 8.400 101.910 10.720 102.120 ;
        RECT 8.560 101.240 10.720 101.910 ;
        RECT 19.770 101.980 20.580 102.250 ;
        RECT 21.390 101.980 22.200 102.790 ;
        RECT 23.280 102.520 23.550 102.790 ;
        RECT 31.700 102.930 33.900 103.430 ;
        RECT 31.700 102.590 34.110 102.930 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 127.360 105.110 129.690 105.430 ;
        RECT 150.750 105.490 152.980 105.690 ;
        RECT 127.360 104.590 129.530 105.110 ;
        RECT 150.750 104.800 152.870 105.490 ;
        RECT 127.180 104.270 129.530 104.590 ;
        RECT 150.620 104.590 152.870 104.800 ;
        RECT 127.180 103.760 129.360 104.270 ;
        RECT 150.620 103.910 152.750 104.590 ;
        RECT 150.480 103.830 152.750 103.910 ;
        RECT 126.980 103.430 129.360 103.760 ;
        RECT 141.420 103.690 152.750 103.830 ;
        RECT 126.980 102.930 129.180 103.430 ;
        RECT 137.430 103.230 139.590 103.500 ;
        RECT 141.420 103.430 152.620 103.690 ;
        RECT 137.430 102.960 139.860 103.230 ;
        RECT 23.280 102.250 23.820 102.520 ;
        RECT 23.010 101.980 23.820 102.250 ;
        RECT 8.560 101.010 10.900 101.240 ;
        RECT 8.720 100.350 10.900 101.010 ;
        RECT 19.770 100.900 23.820 101.980 ;
        RECT 31.900 102.110 34.110 102.590 ;
        RECT 31.900 101.760 34.340 102.110 ;
        RECT 32.110 101.290 34.340 101.760 ;
        RECT 32.110 100.930 34.590 101.290 ;
        RECT 8.720 100.120 11.080 100.350 ;
        RECT 8.900 99.470 11.080 100.120 ;
        RECT 8.900 99.240 11.280 99.470 ;
        RECT 9.080 98.590 11.280 99.240 ;
        RECT 18.620 99.030 19.120 100.720 ;
        RECT 20.040 100.360 23.550 100.900 ;
        RECT 32.340 100.470 34.590 100.930 ;
        RECT 20.580 100.090 23.010 100.360 ;
        RECT 32.340 100.110 34.840 100.470 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 126.770 102.590 129.180 102.930 ;
        RECT 126.770 102.110 128.980 102.590 ;
        RECT 136.890 102.420 140.400 102.960 ;
        RECT 141.420 102.530 141.820 103.430 ;
        RECT 150.480 103.010 152.620 103.430 ;
        RECT 150.320 102.800 152.620 103.010 ;
        RECT 126.540 101.760 128.980 102.110 ;
        RECT 126.540 101.290 128.770 101.760 ;
        RECT 126.290 100.930 128.770 101.290 ;
        RECT 136.620 101.340 140.670 102.420 ;
        RECT 150.320 102.120 152.480 102.800 ;
        RECT 136.620 101.070 137.430 101.340 ;
        RECT 126.290 100.470 128.540 100.930 ;
        RECT 136.620 100.800 137.160 101.070 ;
        RECT 20.850 99.820 23.010 100.090 ;
        RECT 32.590 99.660 34.840 100.110 ;
        RECT 32.590 99.290 35.110 99.660 ;
        RECT 32.840 99.030 35.110 99.290 ;
        RECT 18.620 98.860 35.110 99.030 ;
        RECT 9.080 98.350 11.490 98.590 ;
        RECT 18.620 98.530 35.400 98.860 ;
        RECT 32.840 98.470 35.400 98.530 ;
        RECT 9.280 97.710 11.490 98.350 ;
        RECT 33.110 98.050 35.400 98.470 ;
        RECT 9.280 97.470 11.710 97.710 ;
        RECT 33.110 97.660 35.700 98.050 ;
        RECT 9.490 96.830 11.710 97.470 ;
        RECT 33.400 97.260 35.700 97.660 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
        RECT 126.040 100.110 128.540 100.470 ;
        RECT 136.890 100.530 137.160 100.800 ;
        RECT 138.240 100.530 139.050 101.340 ;
        RECT 139.860 101.070 140.670 101.340 ;
        RECT 150.160 101.910 152.480 102.120 ;
        RECT 150.160 101.240 152.320 101.910 ;
        RECT 140.130 100.800 140.670 101.070 ;
        RECT 149.980 101.010 152.320 101.240 ;
        RECT 140.130 100.530 140.400 100.800 ;
        RECT 136.890 100.260 137.430 100.530 ;
        RECT 137.970 100.260 139.320 100.530 ;
        RECT 139.860 100.260 140.400 100.530 ;
        RECT 149.980 100.350 152.160 101.010 ;
        RECT 126.040 99.660 128.290 100.110 ;
        RECT 137.160 99.990 138.510 100.260 ;
        RECT 138.780 99.990 140.400 100.260 ;
        RECT 149.800 100.120 152.160 100.350 ;
        RECT 137.160 99.720 138.240 99.990 ;
        RECT 139.050 99.720 139.860 99.990 ;
        RECT 125.770 99.290 128.290 99.660 ;
        RECT 125.770 98.860 128.040 99.290 ;
        RECT 137.700 99.180 139.590 99.720 ;
        RECT 149.800 99.470 151.980 100.120 ;
        RECT 149.600 99.240 151.980 99.470 ;
        RECT 136.080 98.910 136.890 99.180 ;
        RECT 137.700 98.910 137.970 99.180 ;
        RECT 138.240 98.910 138.510 99.180 ;
        RECT 138.780 98.910 139.050 99.180 ;
        RECT 139.320 98.910 139.590 99.180 ;
        RECT 140.400 98.910 141.210 99.180 ;
        RECT 125.480 98.470 128.040 98.860 ;
        RECT 125.480 98.050 127.770 98.470 ;
        RECT 135.810 98.370 137.160 98.910 ;
        RECT 140.130 98.370 141.480 98.910 ;
        RECT 149.600 98.590 151.800 99.240 ;
        RECT 136.080 98.100 137.700 98.370 ;
        RECT 139.590 98.100 141.210 98.370 ;
        RECT 149.390 98.350 151.800 98.590 ;
        RECT 125.180 97.660 127.770 98.050 ;
        RECT 136.890 97.830 137.970 98.100 ;
        RECT 139.320 97.830 140.400 98.100 ;
        RECT 33.400 96.860 36.010 97.260 ;
        RECT 9.490 96.590 11.940 96.830 ;
        RECT 9.710 96.310 11.940 96.590 ;
        RECT 33.700 96.470 36.010 96.860 ;
        RECT 9.710 95.910 30.440 96.310 ;
        RECT 33.700 96.050 36.340 96.470 ;
        RECT 9.710 95.710 12.180 95.910 ;
        RECT 9.940 95.090 12.180 95.710 ;
        RECT 9.940 94.830 12.430 95.090 ;
        RECT 10.180 94.230 12.430 94.830 ;
        RECT 26.050 94.880 28.210 95.150 ;
        RECT 26.050 94.610 28.480 94.880 ;
        RECT 10.180 93.960 12.690 94.230 ;
        RECT 25.510 94.070 29.020 94.610 ;
        RECT 30.040 94.180 30.440 95.910 ;
        RECT 34.010 95.680 36.340 96.050 ;
        RECT 34.010 95.260 36.680 95.680 ;
        RECT 34.340 94.910 36.680 95.260 ;
        RECT 34.340 94.470 37.040 94.910 ;
        RECT 34.680 94.130 37.040 94.470 ;
        RECT 10.430 93.370 12.690 93.960 ;
        RECT 10.430 93.090 12.970 93.370 ;
        RECT 10.690 92.510 12.970 93.090 ;
        RECT 25.240 92.990 29.290 94.070 ;
        RECT 34.680 93.680 37.400 94.130 ;
        RECT 25.240 92.720 26.050 92.990 ;
        RECT 10.690 92.230 13.250 92.510 ;
        RECT 25.240 92.450 25.780 92.720 ;
        RECT 10.970 91.650 13.250 92.230 ;
        RECT 25.510 92.180 25.780 92.450 ;
        RECT 26.860 92.180 27.670 92.990 ;
        RECT 28.480 92.720 29.290 92.990 ;
        RECT 35.040 93.370 37.400 93.680 ;
        RECT 35.040 92.910 37.790 93.370 ;
        RECT 28.750 92.450 29.290 92.720 ;
        RECT 35.400 92.610 37.790 92.910 ;
        RECT 28.750 92.180 29.020 92.450 ;
        RECT 25.510 91.910 26.050 92.180 ;
        RECT 26.590 91.910 27.940 92.180 ;
        RECT 28.480 91.910 29.020 92.180 ;
        RECT 35.400 92.130 38.180 92.610 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 125.180 97.260 127.480 97.660 ;
        RECT 137.430 97.560 138.510 97.830 ;
        RECT 138.780 97.560 139.860 97.830 ;
        RECT 149.390 97.710 151.600 98.350 ;
        RECT 124.870 96.860 127.480 97.260 ;
        RECT 137.970 97.020 139.320 97.560 ;
        RECT 149.170 97.470 151.600 97.710 ;
        RECT 124.870 96.470 127.180 96.860 ;
        RECT 137.430 96.750 138.510 97.020 ;
        RECT 138.780 96.750 139.860 97.020 ;
        RECT 149.170 96.830 151.390 97.470 ;
        RECT 124.540 96.050 127.180 96.470 ;
        RECT 135.810 96.480 137.970 96.750 ;
        RECT 139.320 96.480 141.210 96.750 ;
        RECT 148.940 96.590 151.390 96.830 ;
        RECT 135.810 96.210 137.430 96.480 ;
        RECT 139.860 96.210 141.480 96.480 ;
        RECT 124.540 95.680 126.870 96.050 ;
        RECT 124.200 95.260 126.870 95.680 ;
        RECT 135.810 95.940 136.890 96.210 ;
        RECT 140.400 95.940 141.480 96.210 ;
        RECT 148.940 95.960 151.170 96.590 ;
        RECT 135.810 95.670 136.620 95.940 ;
        RECT 140.670 95.670 141.480 95.940 ;
        RECT 148.700 95.710 151.170 95.960 ;
        RECT 136.080 95.400 136.350 95.670 ;
        RECT 137.700 95.400 137.970 95.670 ;
        RECT 138.240 95.400 138.510 95.670 ;
        RECT 138.780 95.400 139.050 95.670 ;
        RECT 139.320 95.400 139.590 95.670 ;
        RECT 140.940 95.400 141.210 95.670 ;
        RECT 124.200 94.910 126.540 95.260 ;
        RECT 123.840 94.470 126.540 94.910 ;
        RECT 137.700 94.860 139.590 95.400 ;
        RECT 148.700 95.090 150.940 95.710 ;
        RECT 137.160 94.590 138.240 94.860 ;
        RECT 139.050 94.590 139.860 94.860 ;
        RECT 148.450 94.830 150.940 95.090 ;
        RECT 123.840 94.130 126.200 94.470 ;
        RECT 137.160 94.320 138.510 94.590 ;
        RECT 138.780 94.320 140.400 94.590 ;
        RECT 123.480 93.680 126.200 94.130 ;
        RECT 136.890 94.050 137.430 94.320 ;
        RECT 137.970 94.050 139.320 94.320 ;
        RECT 139.860 94.050 140.400 94.320 ;
        RECT 148.450 94.230 150.700 94.830 ;
        RECT 136.890 93.780 137.160 94.050 ;
        RECT 123.480 93.370 125.840 93.680 ;
        RECT 123.090 92.910 125.840 93.370 ;
        RECT 136.620 93.510 137.160 93.780 ;
        RECT 136.620 93.240 137.430 93.510 ;
        RECT 138.240 93.240 139.050 94.050 ;
        RECT 140.130 93.780 140.400 94.050 ;
        RECT 148.190 93.960 150.700 94.230 ;
        RECT 140.130 93.510 140.670 93.780 ;
        RECT 139.860 93.240 140.670 93.510 ;
        RECT 148.190 93.370 150.450 93.960 ;
        RECT 123.090 92.610 125.480 92.910 ;
        RECT 10.970 91.370 13.550 91.650 ;
        RECT 25.780 91.640 27.130 91.910 ;
        RECT 27.400 91.640 29.020 91.910 ;
        RECT 35.790 91.860 38.180 92.130 ;
        RECT 25.780 91.370 26.860 91.640 ;
        RECT 27.670 91.370 28.480 91.640 ;
        RECT 35.790 91.370 38.590 91.860 ;
        RECT 11.250 90.800 13.550 91.370 ;
        RECT 26.320 90.830 28.210 91.370 ;
        RECT 36.180 91.110 38.590 91.370 ;
        RECT 11.250 90.510 13.860 90.800 ;
        RECT 24.700 90.560 25.510 90.830 ;
        RECT 26.320 90.560 26.590 90.830 ;
        RECT 26.860 90.560 27.130 90.830 ;
        RECT 27.400 90.560 27.670 90.830 ;
        RECT 27.940 90.560 28.210 90.830 ;
        RECT 29.020 90.560 29.830 90.830 ;
        RECT 36.180 90.610 39.010 91.110 ;
        RECT 11.550 89.950 13.860 90.510 ;
        RECT 24.430 90.020 25.780 90.560 ;
        RECT 28.750 90.020 30.100 90.560 ;
        RECT 36.590 90.380 39.010 90.610 ;
        RECT 11.550 89.650 14.170 89.950 ;
        RECT 24.700 89.750 26.320 90.020 ;
        RECT 28.210 89.750 29.830 90.020 ;
        RECT 36.590 89.860 39.440 90.380 ;
        RECT 11.860 89.110 14.170 89.650 ;
        RECT 25.510 89.480 26.590 89.750 ;
        RECT 27.940 89.480 29.020 89.750 ;
        RECT 37.010 89.650 39.440 89.860 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
        RECT 122.700 92.130 125.480 92.610 ;
        RECT 136.620 92.160 140.670 93.240 ;
        RECT 147.910 93.090 150.450 93.370 ;
        RECT 147.910 92.510 150.190 93.090 ;
        RECT 147.630 92.230 150.190 92.510 ;
        RECT 122.700 91.860 125.090 92.130 ;
        RECT 122.290 91.370 125.090 91.860 ;
        RECT 136.890 91.620 140.400 92.160 ;
        RECT 122.290 91.110 124.700 91.370 ;
        RECT 121.870 90.610 124.700 91.110 ;
        RECT 137.430 91.350 139.860 91.620 ;
        RECT 137.430 91.080 139.590 91.350 ;
        RECT 141.320 91.230 141.820 91.980 ;
        RECT 147.630 91.650 149.910 92.230 ;
        RECT 147.330 91.370 149.910 91.650 ;
        RECT 141.320 90.730 142.600 91.230 ;
        RECT 147.330 90.800 149.630 91.370 ;
        RECT 121.870 90.380 124.290 90.610 ;
        RECT 121.440 90.110 124.290 90.380 ;
        RECT 142.100 90.110 142.600 90.730 ;
        RECT 26.050 89.210 27.130 89.480 ;
        RECT 27.400 89.210 28.480 89.480 ;
        RECT 11.860 88.800 14.500 89.110 ;
        RECT 12.170 88.270 14.500 88.800 ;
        RECT 26.590 88.670 27.940 89.210 ;
        RECT 37.010 89.110 39.890 89.650 ;
        RECT 37.440 88.930 39.890 89.110 ;
        RECT 26.050 88.400 27.130 88.670 ;
        RECT 27.400 88.400 28.480 88.670 ;
        RECT 12.170 87.950 14.840 88.270 ;
        RECT 12.500 87.440 14.840 87.950 ;
        RECT 24.430 88.130 26.590 88.400 ;
        RECT 27.940 88.130 29.830 88.400 ;
        RECT 37.440 88.380 40.350 88.930 ;
        RECT 37.890 88.210 40.350 88.380 ;
        RECT 24.430 87.860 26.050 88.130 ;
        RECT 28.480 87.860 30.100 88.130 ;
        RECT 24.430 87.590 25.510 87.860 ;
        RECT 29.020 87.590 30.100 87.860 ;
        RECT 37.890 87.650 40.820 88.210 ;
        RECT 12.500 87.110 15.190 87.440 ;
        RECT 24.430 87.320 25.240 87.590 ;
        RECT 29.290 87.320 30.100 87.590 ;
        RECT 38.350 87.510 40.820 87.650 ;
        RECT 12.840 86.610 15.190 87.110 ;
        RECT 24.700 87.050 24.970 87.320 ;
        RECT 26.320 87.050 26.590 87.320 ;
        RECT 26.860 87.050 27.130 87.320 ;
        RECT 27.400 87.050 27.670 87.320 ;
        RECT 27.940 87.050 28.210 87.320 ;
        RECT 29.560 87.050 29.830 87.320 ;
        RECT 12.840 86.270 15.550 86.610 ;
        RECT 26.320 86.510 28.210 87.050 ;
        RECT 38.350 86.930 41.310 87.510 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 121.440 89.650 142.600 90.110 ;
        RECT 147.020 90.510 149.630 90.800 ;
        RECT 147.020 89.950 149.330 90.510 ;
        RECT 120.990 89.610 142.600 89.650 ;
        RECT 146.710 89.650 149.330 89.950 ;
        RECT 120.990 89.110 123.870 89.610 ;
        RECT 146.710 89.110 149.020 89.650 ;
        RECT 120.990 88.930 123.440 89.110 ;
        RECT 120.530 88.380 123.440 88.930 ;
        RECT 146.380 88.800 149.020 89.110 ;
        RECT 120.530 88.210 122.990 88.380 ;
        RECT 146.380 88.270 148.710 88.800 ;
        RECT 120.060 87.650 122.990 88.210 ;
        RECT 146.040 87.950 148.710 88.270 ;
        RECT 133.660 87.660 134.060 87.720 ;
        RECT 146.040 87.660 148.380 87.950 ;
        RECT 120.060 87.510 122.530 87.650 ;
        RECT 38.820 86.810 41.310 86.930 ;
        RECT 13.190 85.780 15.550 86.270 ;
        RECT 25.780 86.240 26.860 86.510 ;
        RECT 27.670 86.240 28.480 86.510 ;
        RECT 25.780 85.970 27.130 86.240 ;
        RECT 27.400 85.970 29.020 86.240 ;
        RECT 38.820 86.210 41.800 86.810 ;
        RECT 13.190 85.440 15.920 85.780 ;
        RECT 13.550 84.960 15.920 85.440 ;
        RECT 25.510 85.700 26.050 85.970 ;
        RECT 26.590 85.700 27.940 85.970 ;
        RECT 28.480 85.700 29.020 85.970 ;
        RECT 25.510 85.430 25.780 85.700 ;
        RECT 25.240 85.160 25.780 85.430 ;
        RECT 13.550 84.610 16.300 84.960 ;
        RECT 13.920 84.140 16.300 84.610 ;
        RECT 25.240 84.890 26.050 85.160 ;
        RECT 26.860 84.890 27.670 85.700 ;
        RECT 28.750 85.430 29.020 85.700 ;
        RECT 39.310 86.130 41.800 86.210 ;
        RECT 39.310 85.510 42.310 86.130 ;
        RECT 39.800 85.450 42.310 85.510 ;
        RECT 28.750 85.160 29.290 85.430 ;
        RECT 28.480 84.890 29.290 85.160 ;
        RECT 13.920 83.780 16.690 84.140 ;
        RECT 25.240 83.810 29.290 84.890 ;
        RECT 39.800 84.810 42.830 85.450 ;
        RECT 40.310 84.780 42.830 84.810 ;
        RECT 40.310 84.130 43.360 84.780 ;
        RECT 40.830 84.120 43.360 84.130 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 119.570 86.930 122.530 87.510 ;
        RECT 129.670 87.120 131.830 87.390 ;
        RECT 133.660 87.260 148.380 87.660 ;
        RECT 119.570 86.810 122.060 86.930 ;
        RECT 129.670 86.850 132.100 87.120 ;
        RECT 119.080 86.210 122.060 86.810 ;
        RECT 129.130 86.310 132.640 86.850 ;
        RECT 133.660 86.420 134.060 87.260 ;
        RECT 145.690 87.110 148.380 87.260 ;
        RECT 145.690 86.610 148.040 87.110 ;
        RECT 119.080 86.130 121.570 86.210 ;
        RECT 118.570 85.510 121.570 86.130 ;
        RECT 118.570 85.450 121.080 85.510 ;
        RECT 118.050 84.810 121.080 85.450 ;
        RECT 128.860 85.230 132.910 86.310 ;
        RECT 145.330 86.270 148.040 86.610 ;
        RECT 145.330 85.780 147.690 86.270 ;
        RECT 128.860 84.960 129.670 85.230 ;
        RECT 118.050 84.780 120.570 84.810 ;
        RECT 14.300 83.330 16.690 83.780 ;
        RECT 14.300 82.960 17.090 83.330 ;
        RECT 25.510 83.270 29.020 83.810 ;
        RECT 14.690 82.530 17.090 82.960 ;
        RECT 26.050 83.000 28.480 83.270 ;
        RECT 26.050 82.730 28.210 83.000 ;
        RECT 29.940 82.880 30.440 83.630 ;
        RECT 40.830 83.470 43.910 84.120 ;
        RECT 40.830 83.450 44.460 83.470 ;
        RECT 41.360 82.880 44.460 83.450 ;
        RECT 29.940 82.830 44.460 82.880 ;
        RECT 14.690 82.140 17.500 82.530 ;
        RECT 29.940 82.380 45.030 82.830 ;
        RECT 15.090 81.720 17.500 82.140 ;
        RECT 15.090 81.330 17.920 81.720 ;
        RECT 15.500 80.930 17.920 81.330 ;
        RECT 15.500 80.530 18.350 80.930 ;
        RECT 15.920 80.140 18.350 80.530 ;
        RECT 15.920 79.720 18.790 80.140 ;
        RECT 16.350 79.350 18.790 79.720 ;
        RECT 36.120 79.880 38.280 80.150 ;
        RECT 36.120 79.610 38.550 79.880 ;
        RECT 16.350 78.930 19.240 79.350 ;
        RECT 35.580 79.070 39.090 79.610 ;
        RECT 40.010 79.250 40.510 82.380 ;
        RECT 41.910 82.200 45.030 82.380 ;
        RECT 41.910 82.120 45.610 82.200 ;
        RECT 42.460 81.580 45.610 82.120 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
        RECT 117.520 84.130 120.570 84.780 ;
        RECT 128.860 84.690 129.400 84.960 ;
        RECT 129.130 84.420 129.400 84.690 ;
        RECT 130.480 84.420 131.290 85.230 ;
        RECT 132.100 84.960 132.910 85.230 ;
        RECT 144.960 85.440 147.690 85.780 ;
        RECT 144.960 84.960 147.330 85.440 ;
        RECT 132.370 84.690 132.910 84.960 ;
        RECT 132.370 84.420 132.640 84.690 ;
        RECT 129.130 84.150 129.670 84.420 ;
        RECT 130.210 84.150 131.560 84.420 ;
        RECT 132.100 84.150 132.640 84.420 ;
        RECT 117.520 84.120 120.050 84.130 ;
        RECT 116.970 83.470 120.050 84.120 ;
        RECT 129.400 83.880 130.750 84.150 ;
        RECT 131.020 83.880 132.640 84.150 ;
        RECT 144.580 84.610 147.330 84.960 ;
        RECT 144.580 84.140 146.960 84.610 ;
        RECT 129.400 83.610 130.480 83.880 ;
        RECT 131.290 83.610 132.100 83.880 ;
        RECT 144.190 83.780 146.960 84.140 ;
        RECT 116.420 83.450 120.050 83.470 ;
        RECT 116.420 82.830 119.520 83.450 ;
        RECT 129.940 83.070 131.830 83.610 ;
        RECT 144.190 83.330 146.580 83.780 ;
        RECT 115.850 82.780 119.520 82.830 ;
        RECT 128.320 82.800 129.130 83.070 ;
        RECT 129.940 82.800 130.210 83.070 ;
        RECT 130.480 82.800 130.750 83.070 ;
        RECT 131.020 82.800 131.290 83.070 ;
        RECT 131.560 82.800 131.830 83.070 ;
        RECT 132.640 82.800 133.450 83.070 ;
        RECT 143.790 82.960 146.580 83.330 ;
        RECT 115.850 82.200 118.970 82.780 ;
        RECT 128.050 82.260 129.400 82.800 ;
        RECT 132.370 82.260 133.720 82.800 ;
        RECT 143.790 82.530 146.190 82.960 ;
        RECT 42.460 81.470 46.200 81.580 ;
        RECT 43.030 80.970 46.200 81.470 ;
        RECT 43.030 80.830 46.800 80.970 ;
        RECT 43.610 80.370 46.800 80.830 ;
        RECT 43.610 80.200 47.410 80.370 ;
        RECT 44.200 79.780 47.410 80.200 ;
        RECT 44.200 79.580 48.030 79.780 ;
        RECT 44.800 79.200 48.030 79.580 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 115.270 82.120 118.970 82.200 ;
        RECT 115.270 81.580 118.420 82.120 ;
        RECT 128.320 81.990 129.940 82.260 ;
        RECT 131.830 81.990 133.450 82.260 ;
        RECT 143.380 82.140 146.190 82.530 ;
        RECT 129.130 81.720 130.210 81.990 ;
        RECT 131.560 81.720 132.640 81.990 ;
        RECT 143.380 81.720 145.790 82.140 ;
        RECT 114.680 81.470 118.420 81.580 ;
        RECT 114.680 80.970 117.850 81.470 ;
        RECT 129.670 81.450 130.750 81.720 ;
        RECT 131.020 81.450 132.100 81.720 ;
        RECT 114.080 80.830 117.850 80.970 ;
        RECT 130.210 80.910 131.560 81.450 ;
        RECT 142.960 81.330 145.790 81.720 ;
        RECT 142.960 80.930 145.380 81.330 ;
        RECT 114.080 80.580 117.270 80.830 ;
        RECT 129.670 80.640 130.750 80.910 ;
        RECT 131.020 80.640 132.100 80.910 ;
        RECT 114.080 80.370 127.200 80.580 ;
        RECT 113.470 80.080 127.200 80.370 ;
        RECT 113.470 79.780 116.680 80.080 ;
        RECT 112.850 79.580 116.680 79.780 ;
        RECT 16.790 78.580 19.240 78.930 ;
        RECT 16.790 78.140 19.700 78.580 ;
        RECT 17.240 77.800 19.700 78.140 ;
        RECT 35.310 77.990 39.360 79.070 ;
        RECT 44.800 78.970 48.660 79.200 ;
        RECT 45.410 78.630 48.660 78.970 ;
        RECT 45.410 78.370 49.300 78.630 ;
        RECT 17.240 77.350 20.170 77.800 ;
        RECT 35.310 77.720 36.120 77.990 ;
        RECT 35.310 77.450 35.850 77.720 ;
        RECT 17.700 77.040 20.170 77.350 ;
        RECT 35.580 77.180 35.850 77.450 ;
        RECT 36.930 77.180 37.740 77.990 ;
        RECT 38.550 77.720 39.360 77.990 ;
        RECT 45.630 78.080 49.300 78.370 ;
        RECT 45.630 77.780 49.950 78.080 ;
        RECT 45.630 77.760 46.130 77.780 ;
        RECT 38.820 77.450 39.360 77.720 ;
        RECT 46.660 77.530 49.950 77.780 ;
        RECT 38.820 77.180 39.090 77.450 ;
        RECT 46.660 77.200 50.610 77.530 ;
        RECT 17.700 76.580 20.650 77.040 ;
        RECT 35.580 76.910 36.120 77.180 ;
        RECT 36.660 76.910 38.010 77.180 ;
        RECT 38.550 76.910 39.090 77.180 ;
        RECT 18.170 76.270 20.650 76.580 ;
        RECT 35.850 76.640 37.200 76.910 ;
        RECT 37.470 76.640 39.090 76.910 ;
        RECT 47.300 77.000 50.610 77.200 ;
        RECT 35.850 76.370 36.930 76.640 ;
        RECT 37.740 76.370 38.550 76.640 ;
        RECT 47.300 76.630 51.280 77.000 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
        RECT 112.850 79.200 116.080 79.580 ;
        RECT 112.220 78.970 116.080 79.200 ;
        RECT 112.220 78.630 115.470 78.970 ;
        RECT 111.580 78.370 115.470 78.630 ;
        RECT 111.580 78.080 114.850 78.370 ;
        RECT 110.930 77.780 114.850 78.080 ;
        RECT 110.930 77.530 114.220 77.780 ;
        RECT 110.270 77.200 114.220 77.530 ;
        RECT 110.270 77.000 113.580 77.200 ;
        RECT 47.950 76.480 51.280 76.630 ;
        RECT 109.600 76.630 113.580 77.000 ;
        RECT 109.600 76.480 112.930 76.630 ;
        RECT 18.170 75.800 21.140 76.270 ;
        RECT 36.390 75.830 38.280 76.370 ;
        RECT 47.950 76.080 51.960 76.480 ;
        RECT 48.610 75.970 51.960 76.080 ;
        RECT 108.920 76.080 112.930 76.480 ;
        RECT 108.920 75.970 112.270 76.080 ;
        RECT 18.650 75.520 21.140 75.800 ;
        RECT 34.770 75.560 35.040 75.830 ;
        RECT 36.390 75.560 36.660 75.830 ;
        RECT 36.930 75.560 37.200 75.830 ;
        RECT 37.470 75.560 37.740 75.830 ;
        RECT 38.010 75.560 38.280 75.830 ;
        RECT 39.630 75.560 39.900 75.830 ;
        RECT 18.650 75.040 21.640 75.520 ;
        RECT 19.140 74.770 21.640 75.040 ;
        RECT 34.500 75.290 35.310 75.560 ;
        RECT 39.360 75.290 40.170 75.560 ;
        RECT 48.610 75.530 52.640 75.970 ;
        RECT 34.500 75.020 35.580 75.290 ;
        RECT 39.090 75.020 40.170 75.290 ;
        RECT 19.140 74.270 22.150 74.770 ;
        RECT 34.500 74.750 36.120 75.020 ;
        RECT 38.550 74.750 40.170 75.020 ;
        RECT 49.280 75.480 52.640 75.530 ;
        RECT 108.240 75.530 112.270 75.970 ;
        RECT 108.240 75.480 111.600 75.530 ;
        RECT 49.280 75.000 53.340 75.480 ;
        RECT 49.960 74.990 53.340 75.000 ;
        RECT 107.540 75.000 111.600 75.480 ;
        RECT 107.540 74.990 110.920 75.000 ;
        RECT 34.500 74.480 36.660 74.750 ;
        RECT 38.010 74.480 39.900 74.750 ;
        RECT 49.960 74.520 54.040 74.990 ;
        RECT 106.840 74.520 110.920 74.990 ;
        RECT 49.960 74.480 54.760 74.520 ;
        RECT 19.640 74.030 22.150 74.270 ;
        RECT 36.120 74.210 37.200 74.480 ;
        RECT 37.470 74.210 38.550 74.480 ;
        RECT 19.640 73.520 22.670 74.030 ;
        RECT 36.660 73.670 38.010 74.210 ;
        RECT 50.640 74.060 54.760 74.480 ;
        RECT 106.120 74.480 110.920 74.520 ;
        RECT 106.120 74.060 110.240 74.480 ;
        RECT 50.640 73.970 55.480 74.060 ;
        RECT 20.150 73.290 22.670 73.520 ;
        RECT 36.120 73.400 37.200 73.670 ;
        RECT 37.470 73.400 38.550 73.670 ;
        RECT 51.340 73.610 55.480 73.970 ;
        RECT 105.400 73.970 110.240 74.060 ;
        RECT 105.400 73.610 109.540 73.970 ;
        RECT 51.340 73.480 56.210 73.610 ;
        RECT 20.150 72.770 23.200 73.290 ;
        RECT 35.580 73.130 36.660 73.400 ;
        RECT 38.010 73.130 39.090 73.400 ;
        RECT 52.040 73.180 56.210 73.480 ;
        RECT 104.670 73.480 109.540 73.610 ;
        RECT 117.500 73.790 119.660 74.060 ;
        RECT 117.500 73.520 119.930 73.790 ;
        RECT 104.670 73.180 108.840 73.480 ;
        RECT 34.770 72.860 36.390 73.130 ;
        RECT 38.280 72.860 39.900 73.130 ;
        RECT 52.040 72.990 56.940 73.180 ;
        RECT 20.670 72.570 23.200 72.770 ;
        RECT 20.670 72.030 23.730 72.570 ;
        RECT 34.500 72.320 35.850 72.860 ;
        RECT 38.820 72.320 40.170 72.860 ;
        RECT 52.760 72.760 56.940 72.990 ;
        RECT 103.940 72.990 108.840 73.180 ;
        RECT 103.940 72.760 108.120 72.990 ;
        RECT 116.960 72.980 120.470 73.520 ;
        RECT 121.390 73.160 121.890 80.080 ;
        RECT 126.700 74.250 127.200 80.080 ;
        RECT 128.050 80.370 130.210 80.640 ;
        RECT 131.560 80.370 133.450 80.640 ;
        RECT 142.530 80.530 145.380 80.930 ;
        RECT 128.050 80.100 129.670 80.370 ;
        RECT 132.100 80.100 133.720 80.370 ;
        RECT 142.530 80.140 144.960 80.530 ;
        RECT 128.050 79.830 129.130 80.100 ;
        RECT 132.640 79.830 133.720 80.100 ;
        RECT 128.050 79.560 128.860 79.830 ;
        RECT 132.910 79.560 133.720 79.830 ;
        RECT 142.090 79.720 144.960 80.140 ;
        RECT 128.320 79.290 128.590 79.560 ;
        RECT 129.940 79.290 130.210 79.560 ;
        RECT 130.480 79.290 130.750 79.560 ;
        RECT 131.020 79.290 131.290 79.560 ;
        RECT 131.560 79.290 131.830 79.560 ;
        RECT 133.180 79.290 133.450 79.560 ;
        RECT 142.090 79.350 144.530 79.720 ;
        RECT 129.940 78.750 131.830 79.290 ;
        RECT 141.640 78.930 144.530 79.350 ;
        RECT 129.400 78.480 130.480 78.750 ;
        RECT 131.290 78.480 132.100 78.750 ;
        RECT 141.640 78.580 144.090 78.930 ;
        RECT 129.400 78.210 130.750 78.480 ;
        RECT 131.020 78.210 132.640 78.480 ;
        RECT 129.130 77.940 129.670 78.210 ;
        RECT 130.210 77.940 131.560 78.210 ;
        RECT 132.100 77.940 132.640 78.210 ;
        RECT 129.130 77.670 129.400 77.940 ;
        RECT 128.860 77.400 129.400 77.670 ;
        RECT 128.860 77.130 129.670 77.400 ;
        RECT 130.480 77.130 131.290 77.940 ;
        RECT 132.370 77.670 132.640 77.940 ;
        RECT 141.180 78.140 144.090 78.580 ;
        RECT 141.180 77.800 143.640 78.140 ;
        RECT 132.370 77.400 132.910 77.670 ;
        RECT 132.100 77.130 132.910 77.400 ;
        RECT 128.860 76.050 132.910 77.130 ;
        RECT 140.710 77.350 143.640 77.800 ;
        RECT 140.710 77.040 143.180 77.350 ;
        RECT 140.230 76.580 143.180 77.040 ;
        RECT 140.230 76.270 142.710 76.580 ;
        RECT 129.130 75.510 132.640 76.050 ;
        RECT 129.670 75.240 132.100 75.510 ;
        RECT 129.670 74.970 131.830 75.240 ;
        RECT 133.560 74.250 134.060 75.870 ;
        RECT 139.740 75.800 142.710 76.270 ;
        RECT 139.740 75.520 142.230 75.800 ;
        RECT 139.240 75.040 142.230 75.520 ;
        RECT 139.240 74.770 141.740 75.040 ;
        RECT 126.700 73.750 134.060 74.250 ;
        RECT 138.730 74.270 141.740 74.770 ;
        RECT 138.730 74.030 141.240 74.270 ;
        RECT 138.210 73.520 141.240 74.030 ;
        RECT 138.210 73.290 140.730 73.520 ;
        RECT 52.760 72.520 57.690 72.760 ;
        RECT 53.480 72.350 57.690 72.520 ;
        RECT 103.190 72.520 108.120 72.760 ;
        RECT 103.190 72.350 107.400 72.520 ;
        RECT 34.770 72.050 35.580 72.320 ;
        RECT 36.390 72.050 36.660 72.320 ;
        RECT 36.930 72.050 37.200 72.320 ;
        RECT 37.470 72.050 37.740 72.320 ;
        RECT 38.010 72.050 38.280 72.320 ;
        RECT 39.090 72.050 39.900 72.320 ;
        RECT 53.480 72.060 58.440 72.350 ;
        RECT 21.200 71.840 23.730 72.030 ;
        RECT 21.200 71.290 24.280 71.840 ;
        RECT 36.390 71.510 38.280 72.050 ;
        RECT 53.990 71.960 58.440 72.060 ;
        RECT 102.440 72.060 107.400 72.350 ;
        RECT 102.440 71.960 106.670 72.060 ;
        RECT 53.990 71.610 59.200 71.960 ;
        RECT 21.730 71.130 24.280 71.290 ;
        RECT 35.850 71.240 36.930 71.510 ;
        RECT 37.740 71.240 38.550 71.510 ;
        RECT 21.730 70.570 24.830 71.130 ;
        RECT 35.850 70.970 37.200 71.240 ;
        RECT 37.470 70.970 39.090 71.240 ;
        RECT 22.280 70.420 24.830 70.570 ;
        RECT 35.580 70.700 36.120 70.970 ;
        RECT 36.660 70.700 38.010 70.970 ;
        RECT 38.550 70.700 39.090 70.970 ;
        RECT 35.580 70.430 35.850 70.700 ;
        RECT 22.280 69.840 25.400 70.420 ;
        RECT 22.830 69.720 25.400 69.840 ;
        RECT 35.310 70.160 35.850 70.430 ;
        RECT 35.310 69.890 36.120 70.160 ;
        RECT 36.930 69.890 37.740 70.700 ;
        RECT 38.820 70.430 39.090 70.700 ;
        RECT 38.820 70.160 39.360 70.430 ;
        RECT 38.550 69.890 39.360 70.160 ;
        RECT 22.830 69.130 25.970 69.720 ;
        RECT 23.400 69.030 25.970 69.130 ;
        RECT 23.400 68.420 26.550 69.030 ;
        RECT 35.310 68.810 39.360 69.890 ;
        RECT 23.970 68.340 26.550 68.420 ;
        RECT 23.970 67.720 27.140 68.340 ;
        RECT 35.580 68.270 39.090 68.810 ;
        RECT 50.100 68.730 52.260 69.000 ;
        RECT 36.120 68.000 38.550 68.270 ;
        RECT 36.120 67.730 38.280 68.000 ;
        RECT 24.550 67.660 27.140 67.720 ;
        RECT 24.550 67.030 27.740 67.660 ;
        RECT 25.140 66.990 27.740 67.030 ;
        RECT 25.140 66.340 28.340 66.990 ;
        RECT 25.740 66.330 28.340 66.340 ;
        RECT 25.740 65.670 28.960 66.330 ;
        RECT 25.740 65.660 29.580 65.670 ;
        RECT 26.340 65.020 29.580 65.660 ;
        RECT 26.340 64.990 30.210 65.020 ;
        RECT 26.960 64.380 30.210 64.990 ;
        RECT 26.960 64.330 30.850 64.380 ;
        RECT 27.580 63.750 30.850 64.330 ;
        RECT 27.580 63.670 31.500 63.750 ;
        RECT 28.210 63.130 31.500 63.670 ;
        RECT 28.210 63.020 32.160 63.130 ;
        RECT 28.850 62.510 32.160 63.020 ;
        RECT 28.850 62.380 32.820 62.510 ;
        RECT 29.500 61.910 32.820 62.380 ;
        RECT 29.500 61.750 33.490 61.910 ;
        RECT 30.160 61.310 33.490 61.750 ;
        RECT 30.160 61.130 34.170 61.310 ;
        RECT 30.820 60.720 34.170 61.130 ;
        RECT 30.820 60.510 34.860 60.720 ;
        RECT 31.490 60.140 34.860 60.510 ;
        RECT 31.490 59.910 35.550 60.140 ;
        RECT 32.170 59.570 35.550 59.910 ;
        RECT 32.170 59.310 36.250 59.570 ;
        RECT 32.860 59.000 36.250 59.310 ;
        RECT 32.860 58.720 36.960 59.000 ;
        RECT 33.550 58.450 36.960 58.720 ;
        RECT 33.550 58.140 37.670 58.450 ;
        RECT 34.250 57.900 37.670 58.140 ;
        RECT 34.250 57.570 38.400 57.900 ;
        RECT 34.960 57.370 38.400 57.570 ;
        RECT 34.960 57.000 39.120 57.370 ;
        RECT 35.670 56.840 39.120 57.000 ;
        RECT 35.670 56.450 39.860 56.840 ;
        RECT 36.400 56.320 39.860 56.450 ;
        RECT 40.110 56.320 40.510 68.700 ;
        RECT 50.100 68.460 52.530 68.730 ;
        RECT 49.560 67.920 53.070 68.460 ;
        RECT 53.990 68.100 54.490 71.610 ;
        RECT 54.940 71.570 59.200 71.610 ;
        RECT 101.680 71.610 106.670 71.960 ;
        RECT 116.690 71.900 120.740 72.980 ;
        RECT 137.680 72.770 140.730 73.290 ;
        RECT 137.680 72.570 140.210 72.770 ;
        RECT 116.690 71.630 117.500 71.900 ;
        RECT 101.680 71.570 106.410 71.610 ;
        RECT 54.940 71.210 59.960 71.570 ;
        RECT 100.920 71.210 106.410 71.570 ;
        RECT 116.690 71.360 117.230 71.630 ;
        RECT 54.940 71.180 60.740 71.210 ;
        RECT 55.690 70.850 60.740 71.180 ;
        RECT 100.140 71.180 106.410 71.210 ;
        RECT 100.140 70.850 105.190 71.180 ;
        RECT 55.690 70.760 61.510 70.850 ;
        RECT 56.440 70.510 61.510 70.760 ;
        RECT 99.370 70.760 105.190 70.850 ;
        RECT 99.370 70.510 104.440 70.760 ;
        RECT 56.440 70.350 62.300 70.510 ;
        RECT 57.200 70.180 62.300 70.350 ;
        RECT 98.580 70.350 104.440 70.510 ;
        RECT 98.580 70.180 103.680 70.350 ;
        RECT 57.200 69.960 63.090 70.180 ;
        RECT 57.960 69.870 63.090 69.960 ;
        RECT 97.790 69.960 103.680 70.180 ;
        RECT 97.790 69.870 102.920 69.960 ;
        RECT 57.960 69.570 63.880 69.870 ;
        RECT 97.000 69.570 102.920 69.870 ;
        RECT 58.740 69.280 64.690 69.570 ;
        RECT 96.190 69.280 102.140 69.570 ;
        RECT 58.740 69.210 65.490 69.280 ;
        RECT 59.510 69.010 65.490 69.210 ;
        RECT 95.390 69.210 102.140 69.280 ;
        RECT 95.390 69.010 101.370 69.210 ;
        RECT 59.510 68.850 66.300 69.010 ;
        RECT 60.300 68.760 66.300 68.850 ;
        RECT 94.580 68.850 101.370 69.010 ;
        RECT 94.580 68.760 100.580 68.850 ;
        RECT 60.300 68.510 67.120 68.760 ;
        RECT 93.760 68.510 100.580 68.760 ;
        RECT 61.090 68.280 67.940 68.510 ;
        RECT 92.940 68.280 99.790 68.510 ;
        RECT 61.090 68.180 68.760 68.280 ;
        RECT 61.880 68.070 68.760 68.180 ;
        RECT 92.120 68.180 99.790 68.280 ;
        RECT 92.120 68.070 99.000 68.180 ;
        RECT 49.290 66.840 53.340 67.920 ;
        RECT 61.880 67.870 69.590 68.070 ;
        RECT 91.290 67.870 99.000 68.070 ;
        RECT 62.690 67.690 70.420 67.870 ;
        RECT 90.460 67.690 98.190 67.870 ;
        RECT 62.690 67.570 71.260 67.690 ;
        RECT 63.490 67.520 71.260 67.570 ;
        RECT 89.620 67.570 98.190 67.690 ;
        RECT 89.620 67.520 97.390 67.570 ;
        RECT 63.490 67.360 72.100 67.520 ;
        RECT 88.780 67.360 97.390 67.520 ;
        RECT 63.490 67.280 72.940 67.360 ;
        RECT 64.300 67.220 72.940 67.280 ;
        RECT 87.940 67.280 97.390 67.360 ;
        RECT 87.940 67.220 96.580 67.280 ;
        RECT 64.300 67.090 73.780 67.220 ;
        RECT 87.100 67.090 96.580 67.220 ;
        RECT 64.300 67.010 74.630 67.090 ;
        RECT 49.290 66.570 50.100 66.840 ;
        RECT 49.290 66.300 49.830 66.570 ;
        RECT 49.560 66.030 49.830 66.300 ;
        RECT 50.910 66.030 51.720 66.840 ;
        RECT 52.530 66.570 53.340 66.840 ;
        RECT 65.120 66.980 74.630 67.010 ;
        RECT 86.250 67.010 96.580 67.090 ;
        RECT 86.250 66.980 95.760 67.010 ;
        RECT 65.120 66.880 75.470 66.980 ;
        RECT 85.410 66.880 95.760 66.980 ;
        RECT 65.120 66.800 76.320 66.880 ;
        RECT 84.560 66.800 95.760 66.880 ;
        RECT 65.120 66.760 77.170 66.800 ;
        RECT 52.800 66.300 53.340 66.570 ;
        RECT 65.940 66.730 77.170 66.760 ;
        RECT 83.710 66.760 95.760 66.800 ;
        RECT 83.710 66.730 94.940 66.760 ;
        RECT 65.940 66.680 78.030 66.730 ;
        RECT 82.850 66.680 94.940 66.730 ;
        RECT 65.940 66.640 78.880 66.680 ;
        RECT 82.000 66.640 94.940 66.680 ;
        RECT 65.940 66.620 79.730 66.640 ;
        RECT 81.150 66.620 94.940 66.640 ;
        RECT 65.940 66.510 94.940 66.620 ;
        RECT 52.800 66.030 53.070 66.300 ;
        RECT 66.760 66.280 94.120 66.510 ;
        RECT 67.590 66.070 93.290 66.280 ;
        RECT 49.560 65.760 50.100 66.030 ;
        RECT 50.640 65.760 51.990 66.030 ;
        RECT 52.530 65.760 53.070 66.030 ;
        RECT 68.420 65.870 92.460 66.070 ;
        RECT 49.830 65.490 51.180 65.760 ;
        RECT 51.450 65.490 53.070 65.760 ;
        RECT 69.260 65.690 91.620 65.870 ;
        RECT 70.100 65.520 90.780 65.690 ;
        RECT 49.830 65.220 50.910 65.490 ;
        RECT 51.720 65.220 52.530 65.490 ;
        RECT 70.640 65.360 89.940 65.520 ;
        RECT 50.370 64.680 52.260 65.220 ;
        RECT 48.750 64.410 49.020 64.680 ;
        RECT 50.370 64.410 50.640 64.680 ;
        RECT 50.910 64.410 51.180 64.680 ;
        RECT 51.450 64.410 51.720 64.680 ;
        RECT 51.990 64.410 52.260 64.680 ;
        RECT 53.610 64.410 53.880 64.680 ;
        RECT 48.480 64.140 49.290 64.410 ;
        RECT 53.340 64.140 54.150 64.410 ;
        RECT 48.480 63.870 49.560 64.140 ;
        RECT 53.070 63.870 54.150 64.140 ;
        RECT 48.480 63.600 50.100 63.870 ;
        RECT 52.530 63.600 54.150 63.870 ;
        RECT 48.480 63.330 50.640 63.600 ;
        RECT 51.990 63.330 53.880 63.600 ;
        RECT 50.100 63.060 51.180 63.330 ;
        RECT 51.450 63.060 52.530 63.330 ;
        RECT 50.640 62.520 51.990 63.060 ;
        RECT 50.100 62.250 51.180 62.520 ;
        RECT 51.450 62.250 52.530 62.520 ;
        RECT 49.560 61.980 50.640 62.250 ;
        RECT 51.990 61.980 53.070 62.250 ;
        RECT 66.750 62.200 68.910 62.470 ;
        RECT 48.750 61.710 50.370 61.980 ;
        RECT 52.260 61.710 53.880 61.980 ;
        RECT 66.750 61.930 69.180 62.200 ;
        RECT 48.480 61.170 49.830 61.710 ;
        RECT 52.800 61.170 54.150 61.710 ;
        RECT 66.210 61.390 69.720 61.930 ;
        RECT 70.640 61.570 71.140 65.360 ;
        RECT 71.780 65.220 89.100 65.360 ;
        RECT 72.630 65.090 88.250 65.220 ;
        RECT 73.470 64.980 87.410 65.090 ;
        RECT 74.320 64.880 86.560 64.980 ;
        RECT 75.170 64.800 85.710 64.880 ;
        RECT 76.030 64.730 84.850 64.800 ;
        RECT 76.880 64.680 84.000 64.730 ;
        RECT 77.730 64.640 83.150 64.680 ;
        RECT 78.590 64.620 82.290 64.640 ;
        RECT 79.440 64.610 81.430 64.620 ;
        RECT 48.750 60.900 49.560 61.170 ;
        RECT 50.370 60.900 50.640 61.170 ;
        RECT 50.910 60.900 51.180 61.170 ;
        RECT 51.450 60.900 51.720 61.170 ;
        RECT 51.990 60.900 52.260 61.170 ;
        RECT 53.070 60.900 53.880 61.170 ;
        RECT 50.370 60.360 52.260 60.900 ;
        RECT 49.830 60.090 50.910 60.360 ;
        RECT 51.720 60.090 52.530 60.360 ;
        RECT 65.940 60.310 69.990 61.390 ;
        RECT 84.580 60.860 86.740 61.130 ;
        RECT 84.580 60.590 87.010 60.860 ;
        RECT 49.830 59.820 51.180 60.090 ;
        RECT 51.450 59.820 53.070 60.090 ;
        RECT 49.560 59.550 50.100 59.820 ;
        RECT 50.640 59.550 51.990 59.820 ;
        RECT 52.530 59.550 53.070 59.820 ;
        RECT 65.940 60.040 66.750 60.310 ;
        RECT 65.940 59.770 66.480 60.040 ;
        RECT 49.560 59.280 49.830 59.550 ;
        RECT 49.290 59.010 49.830 59.280 ;
        RECT 49.290 58.740 50.100 59.010 ;
        RECT 50.910 58.740 51.720 59.550 ;
        RECT 52.800 59.280 53.070 59.550 ;
        RECT 66.210 59.500 66.480 59.770 ;
        RECT 67.560 59.500 68.370 60.310 ;
        RECT 69.180 60.040 69.990 60.310 ;
        RECT 84.040 60.050 87.550 60.590 ;
        RECT 88.470 60.230 88.970 65.220 ;
        RECT 102.020 64.840 104.180 65.110 ;
        RECT 102.020 64.570 104.450 64.840 ;
        RECT 101.480 64.030 104.990 64.570 ;
        RECT 105.910 64.210 106.410 71.180 ;
        RECT 116.960 71.090 117.230 71.360 ;
        RECT 118.310 71.090 119.120 71.900 ;
        RECT 119.930 71.630 120.740 71.900 ;
        RECT 137.150 72.030 140.210 72.570 ;
        RECT 137.150 71.840 139.680 72.030 ;
        RECT 120.200 71.360 120.740 71.630 ;
        RECT 120.200 71.090 120.470 71.360 ;
        RECT 136.600 71.290 139.680 71.840 ;
        RECT 136.600 71.130 139.150 71.290 ;
        RECT 116.960 70.820 117.500 71.090 ;
        RECT 118.040 70.820 119.390 71.090 ;
        RECT 119.930 70.820 120.470 71.090 ;
        RECT 117.230 70.550 118.580 70.820 ;
        RECT 118.850 70.550 120.470 70.820 ;
        RECT 136.050 70.570 139.150 71.130 ;
        RECT 117.230 70.280 118.310 70.550 ;
        RECT 119.120 70.280 119.930 70.550 ;
        RECT 136.050 70.420 138.600 70.570 ;
        RECT 117.770 69.740 119.660 70.280 ;
        RECT 135.480 69.840 138.600 70.420 ;
        RECT 116.150 69.470 116.420 69.740 ;
        RECT 117.770 69.470 118.040 69.740 ;
        RECT 118.310 69.470 118.580 69.740 ;
        RECT 118.850 69.470 119.120 69.740 ;
        RECT 119.390 69.470 119.660 69.740 ;
        RECT 121.010 69.470 121.280 69.740 ;
        RECT 135.480 69.720 138.050 69.840 ;
        RECT 115.880 69.200 116.690 69.470 ;
        RECT 120.740 69.200 121.550 69.470 ;
        RECT 115.880 68.930 116.960 69.200 ;
        RECT 120.470 68.930 121.550 69.200 ;
        RECT 134.910 69.130 138.050 69.720 ;
        RECT 134.910 69.030 137.480 69.130 ;
        RECT 115.880 68.660 117.500 68.930 ;
        RECT 119.930 68.660 121.550 68.930 ;
        RECT 115.880 68.390 118.040 68.660 ;
        RECT 119.390 68.390 121.280 68.660 ;
        RECT 134.330 68.420 137.480 69.030 ;
        RECT 117.500 68.120 118.580 68.390 ;
        RECT 118.850 68.120 119.930 68.390 ;
        RECT 134.330 68.340 136.910 68.420 ;
        RECT 118.040 67.580 119.390 68.120 ;
        RECT 133.740 67.720 136.910 68.340 ;
        RECT 133.740 67.660 136.330 67.720 ;
        RECT 117.500 67.310 118.580 67.580 ;
        RECT 118.850 67.310 119.930 67.580 ;
        RECT 116.960 67.040 118.040 67.310 ;
        RECT 119.390 67.040 120.470 67.310 ;
        RECT 116.150 66.770 117.770 67.040 ;
        RECT 119.660 66.770 121.280 67.040 ;
        RECT 133.140 67.030 136.330 67.660 ;
        RECT 133.140 66.990 135.740 67.030 ;
        RECT 115.880 66.230 117.230 66.770 ;
        RECT 120.200 66.230 121.550 66.770 ;
        RECT 132.540 66.340 135.740 66.990 ;
        RECT 132.540 66.330 135.140 66.340 ;
        RECT 116.150 65.960 116.960 66.230 ;
        RECT 117.770 65.960 118.040 66.230 ;
        RECT 118.310 65.960 118.580 66.230 ;
        RECT 118.850 65.960 119.120 66.230 ;
        RECT 119.390 65.960 119.660 66.230 ;
        RECT 120.470 65.960 121.280 66.230 ;
        RECT 117.770 65.420 119.660 65.960 ;
        RECT 131.920 65.670 135.140 66.330 ;
        RECT 131.300 65.660 135.140 65.670 ;
        RECT 117.230 65.150 118.310 65.420 ;
        RECT 119.120 65.150 119.930 65.420 ;
        RECT 117.230 64.880 118.580 65.150 ;
        RECT 118.850 64.880 120.470 65.150 ;
        RECT 131.300 65.020 134.540 65.660 ;
        RECT 116.960 64.610 117.500 64.880 ;
        RECT 118.040 64.610 119.390 64.880 ;
        RECT 119.930 64.610 120.470 64.880 ;
        RECT 116.960 64.340 117.230 64.610 ;
        RECT 116.690 64.070 117.230 64.340 ;
        RECT 101.210 62.950 105.260 64.030 ;
        RECT 101.210 62.680 102.020 62.950 ;
        RECT 101.210 62.410 101.750 62.680 ;
        RECT 101.480 62.140 101.750 62.410 ;
        RECT 102.830 62.140 103.640 62.950 ;
        RECT 104.450 62.680 105.260 62.950 ;
        RECT 116.690 63.800 117.500 64.070 ;
        RECT 118.310 63.800 119.120 64.610 ;
        RECT 120.200 64.340 120.470 64.610 ;
        RECT 130.670 64.990 134.540 65.020 ;
        RECT 130.670 64.380 133.920 64.990 ;
        RECT 120.200 64.070 120.740 64.340 ;
        RECT 119.930 63.800 120.740 64.070 ;
        RECT 116.690 62.720 120.740 63.800 ;
        RECT 130.030 64.330 133.920 64.380 ;
        RECT 130.030 63.750 133.300 64.330 ;
        RECT 129.380 63.670 133.300 63.750 ;
        RECT 129.380 63.130 132.670 63.670 ;
        RECT 128.720 63.020 132.670 63.130 ;
        RECT 104.720 62.410 105.260 62.680 ;
        RECT 104.720 62.140 104.990 62.410 ;
        RECT 116.960 62.180 120.470 62.720 ;
        RECT 101.480 61.870 102.020 62.140 ;
        RECT 102.560 61.870 103.910 62.140 ;
        RECT 104.450 61.870 104.990 62.140 ;
        RECT 101.750 61.600 103.100 61.870 ;
        RECT 103.370 61.600 104.990 61.870 ;
        RECT 117.500 61.910 119.930 62.180 ;
        RECT 117.500 61.640 119.660 61.910 ;
        RECT 101.750 61.330 102.830 61.600 ;
        RECT 103.640 61.330 104.450 61.600 ;
        RECT 102.290 60.790 104.180 61.330 ;
        RECT 100.670 60.520 100.940 60.790 ;
        RECT 102.290 60.520 102.560 60.790 ;
        RECT 102.830 60.520 103.100 60.790 ;
        RECT 103.370 60.520 103.640 60.790 ;
        RECT 103.910 60.520 104.180 60.790 ;
        RECT 105.530 60.520 105.800 60.790 ;
        RECT 100.400 60.250 101.210 60.520 ;
        RECT 105.260 60.250 106.070 60.520 ;
        RECT 69.450 59.770 69.990 60.040 ;
        RECT 69.450 59.500 69.720 59.770 ;
        RECT 52.800 59.010 53.340 59.280 ;
        RECT 66.210 59.230 66.750 59.500 ;
        RECT 67.290 59.230 68.640 59.500 ;
        RECT 69.180 59.230 69.720 59.500 ;
        RECT 52.530 58.740 53.340 59.010 ;
        RECT 49.290 57.660 53.340 58.740 ;
        RECT 66.480 58.960 67.830 59.230 ;
        RECT 68.100 58.960 69.720 59.230 ;
        RECT 83.770 58.970 87.820 60.050 ;
        RECT 100.400 59.980 101.480 60.250 ;
        RECT 104.990 59.980 106.070 60.250 ;
        RECT 100.400 59.710 102.020 59.980 ;
        RECT 104.450 59.710 106.070 59.980 ;
        RECT 100.400 59.440 102.560 59.710 ;
        RECT 103.910 59.440 105.800 59.710 ;
        RECT 102.020 59.170 103.100 59.440 ;
        RECT 103.370 59.170 104.450 59.440 ;
        RECT 66.480 58.690 67.560 58.960 ;
        RECT 68.370 58.690 69.180 58.960 ;
        RECT 83.770 58.700 84.580 58.970 ;
        RECT 67.020 58.150 68.910 58.690 ;
        RECT 83.770 58.430 84.310 58.700 ;
        RECT 84.040 58.160 84.310 58.430 ;
        RECT 85.390 58.160 86.200 58.970 ;
        RECT 87.010 58.700 87.820 58.970 ;
        RECT 87.280 58.430 87.820 58.700 ;
        RECT 102.560 58.630 103.910 59.170 ;
        RECT 87.280 58.160 87.550 58.430 ;
        RECT 102.020 58.360 103.100 58.630 ;
        RECT 103.370 58.360 104.450 58.630 ;
        RECT 65.400 57.880 65.670 58.150 ;
        RECT 67.020 57.880 67.290 58.150 ;
        RECT 67.560 57.880 67.830 58.150 ;
        RECT 68.100 57.880 68.370 58.150 ;
        RECT 68.640 57.880 68.910 58.150 ;
        RECT 70.260 57.880 70.530 58.150 ;
        RECT 84.040 57.890 84.580 58.160 ;
        RECT 85.120 57.890 86.470 58.160 ;
        RECT 87.010 57.890 87.550 58.160 ;
        RECT 101.480 58.090 102.560 58.360 ;
        RECT 103.910 58.090 104.990 58.360 ;
        RECT 49.560 57.120 53.070 57.660 ;
        RECT 65.130 57.610 65.940 57.880 ;
        RECT 69.990 57.610 70.800 57.880 ;
        RECT 50.100 56.850 52.530 57.120 ;
        RECT 50.100 56.580 52.260 56.850 ;
        RECT 36.400 55.900 40.600 56.320 ;
        RECT 37.120 55.810 40.600 55.900 ;
        RECT 37.120 55.370 41.350 55.810 ;
        RECT 37.860 55.310 41.350 55.370 ;
        RECT 37.860 54.840 42.100 55.310 ;
        RECT 38.600 54.820 42.100 54.840 ;
        RECT 38.600 54.340 42.870 54.820 ;
        RECT 38.600 54.320 43.630 54.340 ;
        RECT 39.350 53.870 43.630 54.320 ;
        RECT 39.350 53.810 44.410 53.870 ;
        RECT 40.100 53.410 44.410 53.810 ;
        RECT 40.100 53.310 45.180 53.410 ;
        RECT 40.870 52.960 45.180 53.310 ;
        RECT 40.870 52.820 45.970 52.960 ;
        RECT 41.630 52.520 45.970 52.820 ;
        RECT 41.630 52.340 46.760 52.520 ;
        RECT 42.410 52.090 46.760 52.340 ;
        RECT 42.410 51.870 47.550 52.090 ;
        RECT 43.180 51.670 47.550 51.870 ;
        RECT 43.180 51.410 48.360 51.670 ;
        RECT 43.970 51.260 48.360 51.410 ;
        RECT 43.970 50.960 49.160 51.260 ;
        RECT 44.760 50.860 49.160 50.960 ;
        RECT 44.760 50.520 49.970 50.860 ;
        RECT 45.550 50.470 49.970 50.520 ;
        RECT 45.550 50.090 50.790 50.470 ;
        RECT 46.360 49.720 51.610 50.090 ;
        RECT 46.360 49.670 52.440 49.720 ;
        RECT 47.160 49.360 52.440 49.670 ;
        RECT 47.160 49.260 53.270 49.360 ;
        RECT 47.970 49.010 53.270 49.260 ;
        RECT 54.090 49.010 54.490 57.550 ;
        RECT 65.130 57.340 66.210 57.610 ;
        RECT 69.720 57.340 70.800 57.610 ;
        RECT 84.310 57.620 85.660 57.890 ;
        RECT 85.930 57.620 87.550 57.890 ;
        RECT 100.670 57.820 102.290 58.090 ;
        RECT 104.180 57.820 105.800 58.090 ;
        RECT 84.310 57.350 85.390 57.620 ;
        RECT 86.200 57.350 87.010 57.620 ;
        RECT 65.130 57.070 66.750 57.340 ;
        RECT 69.180 57.070 70.800 57.340 ;
        RECT 65.130 56.800 67.290 57.070 ;
        RECT 68.640 56.800 70.530 57.070 ;
        RECT 84.850 56.810 86.740 57.350 ;
        RECT 100.400 57.280 101.750 57.820 ;
        RECT 104.720 57.280 106.070 57.820 ;
        RECT 121.490 57.370 121.890 62.610 ;
        RECT 128.720 62.510 132.030 63.020 ;
        RECT 128.060 62.380 132.030 62.510 ;
        RECT 128.060 61.910 131.380 62.380 ;
        RECT 127.390 61.750 131.380 61.910 ;
        RECT 127.390 61.310 130.720 61.750 ;
        RECT 126.710 61.130 130.720 61.310 ;
        RECT 126.710 60.720 130.060 61.130 ;
        RECT 126.020 60.510 130.060 60.720 ;
        RECT 126.020 60.140 129.390 60.510 ;
        RECT 125.330 59.910 129.390 60.140 ;
        RECT 125.330 59.570 128.710 59.910 ;
        RECT 124.630 59.310 128.710 59.570 ;
        RECT 124.630 59.000 128.020 59.310 ;
        RECT 123.920 58.720 128.020 59.000 ;
        RECT 123.920 58.450 127.330 58.720 ;
        RECT 123.210 58.140 127.330 58.450 ;
        RECT 123.210 57.900 126.630 58.140 ;
        RECT 122.480 57.570 126.630 57.900 ;
        RECT 122.480 57.370 125.920 57.570 ;
        RECT 100.670 57.010 101.480 57.280 ;
        RECT 102.290 57.010 102.560 57.280 ;
        RECT 102.830 57.010 103.100 57.280 ;
        RECT 103.370 57.010 103.640 57.280 ;
        RECT 103.910 57.010 104.180 57.280 ;
        RECT 104.990 57.010 105.800 57.280 ;
        RECT 66.750 56.530 67.830 56.800 ;
        RECT 68.100 56.530 69.180 56.800 ;
        RECT 83.230 56.540 83.500 56.810 ;
        RECT 84.850 56.540 85.120 56.810 ;
        RECT 85.390 56.540 85.660 56.810 ;
        RECT 85.930 56.540 86.200 56.810 ;
        RECT 86.470 56.540 86.740 56.810 ;
        RECT 88.090 56.540 88.360 56.810 ;
        RECT 67.290 55.990 68.640 56.530 ;
        RECT 82.960 56.270 83.770 56.540 ;
        RECT 87.820 56.270 88.630 56.540 ;
        RECT 102.290 56.470 104.180 57.010 ;
        RECT 121.490 57.000 125.920 57.370 ;
        RECT 121.490 56.840 125.210 57.000 ;
        RECT 82.960 56.000 84.040 56.270 ;
        RECT 87.550 56.000 88.630 56.270 ;
        RECT 66.750 55.720 67.830 55.990 ;
        RECT 68.100 55.720 69.180 55.990 ;
        RECT 82.960 55.730 84.580 56.000 ;
        RECT 87.010 55.730 88.630 56.000 ;
        RECT 101.750 56.200 102.830 56.470 ;
        RECT 103.640 56.200 104.450 56.470 ;
        RECT 121.020 56.450 125.210 56.840 ;
        RECT 121.020 56.320 124.480 56.450 ;
        RECT 101.750 55.930 103.100 56.200 ;
        RECT 103.370 55.930 104.990 56.200 ;
        RECT 66.210 55.450 67.290 55.720 ;
        RECT 68.640 55.450 69.720 55.720 ;
        RECT 82.960 55.460 85.120 55.730 ;
        RECT 86.470 55.460 88.360 55.730 ;
        RECT 101.480 55.660 102.020 55.930 ;
        RECT 102.560 55.660 103.910 55.930 ;
        RECT 104.450 55.660 104.990 55.930 ;
        RECT 120.280 55.900 124.480 56.320 ;
        RECT 120.280 55.810 123.760 55.900 ;
        RECT 65.400 55.180 67.020 55.450 ;
        RECT 68.910 55.180 70.530 55.450 ;
        RECT 84.580 55.190 85.660 55.460 ;
        RECT 85.930 55.190 87.010 55.460 ;
        RECT 101.480 55.390 101.750 55.660 ;
        RECT 65.130 54.640 66.480 55.180 ;
        RECT 69.450 54.640 70.800 55.180 ;
        RECT 85.120 54.650 86.470 55.190 ;
        RECT 101.210 55.120 101.750 55.390 ;
        RECT 101.210 54.850 102.020 55.120 ;
        RECT 102.830 54.850 103.640 55.660 ;
        RECT 104.720 55.390 104.990 55.660 ;
        RECT 104.720 55.120 105.260 55.390 ;
        RECT 119.530 55.370 123.760 55.810 ;
        RECT 119.530 55.310 123.020 55.370 ;
        RECT 104.450 54.850 105.260 55.120 ;
        RECT 65.400 54.370 66.210 54.640 ;
        RECT 67.020 54.370 67.290 54.640 ;
        RECT 67.560 54.370 67.830 54.640 ;
        RECT 68.100 54.370 68.370 54.640 ;
        RECT 68.640 54.370 68.910 54.640 ;
        RECT 69.720 54.370 70.530 54.640 ;
        RECT 84.580 54.380 85.660 54.650 ;
        RECT 85.930 54.380 87.010 54.650 ;
        RECT 67.020 53.830 68.910 54.370 ;
        RECT 84.040 54.110 85.120 54.380 ;
        RECT 86.470 54.110 87.550 54.380 ;
        RECT 83.230 53.840 84.850 54.110 ;
        RECT 86.740 53.840 88.360 54.110 ;
        RECT 66.480 53.560 67.560 53.830 ;
        RECT 68.370 53.560 69.180 53.830 ;
        RECT 66.480 53.290 67.830 53.560 ;
        RECT 68.100 53.290 69.720 53.560 ;
        RECT 82.960 53.300 84.310 53.840 ;
        RECT 87.280 53.300 88.630 53.840 ;
        RECT 101.210 53.770 105.260 54.850 ;
        RECT 118.780 54.840 123.020 55.310 ;
        RECT 118.780 54.820 122.280 54.840 ;
        RECT 118.010 54.340 122.280 54.820 ;
        RECT 117.250 54.320 122.280 54.340 ;
        RECT 117.250 53.870 121.530 54.320 ;
        RECT 116.470 53.810 121.530 53.870 ;
        RECT 66.210 53.020 66.750 53.290 ;
        RECT 67.290 53.020 68.640 53.290 ;
        RECT 69.180 53.020 69.720 53.290 ;
        RECT 83.230 53.030 84.040 53.300 ;
        RECT 84.850 53.030 85.120 53.300 ;
        RECT 85.390 53.030 85.660 53.300 ;
        RECT 85.930 53.030 86.200 53.300 ;
        RECT 86.470 53.030 86.740 53.300 ;
        RECT 87.550 53.030 88.360 53.300 ;
        RECT 101.480 53.230 104.990 53.770 ;
        RECT 66.210 52.750 66.480 53.020 ;
        RECT 65.940 52.480 66.480 52.750 ;
        RECT 65.940 52.210 66.750 52.480 ;
        RECT 67.560 52.210 68.370 53.020 ;
        RECT 69.450 52.750 69.720 53.020 ;
        RECT 69.450 52.480 69.990 52.750 ;
        RECT 84.850 52.490 86.740 53.030 ;
        RECT 102.020 52.960 104.450 53.230 ;
        RECT 102.020 52.690 104.180 52.960 ;
        RECT 69.180 52.210 69.990 52.480 ;
        RECT 65.940 51.130 69.990 52.210 ;
        RECT 84.310 52.220 85.390 52.490 ;
        RECT 86.200 52.220 87.010 52.490 ;
        RECT 84.310 51.950 85.660 52.220 ;
        RECT 85.930 51.950 87.550 52.220 ;
        RECT 84.040 51.680 84.580 51.950 ;
        RECT 85.120 51.680 86.470 51.950 ;
        RECT 87.010 51.680 87.550 51.950 ;
        RECT 84.040 51.410 84.310 51.680 ;
        RECT 83.770 51.140 84.310 51.410 ;
        RECT 66.210 50.590 69.720 51.130 ;
        RECT 66.750 50.320 69.180 50.590 ;
        RECT 66.750 50.050 68.910 50.320 ;
        RECT 47.970 48.860 54.490 49.010 ;
        RECT 48.790 48.670 54.490 48.860 ;
        RECT 48.790 48.470 54.940 48.670 ;
        RECT 49.610 48.340 54.940 48.470 ;
        RECT 49.610 48.090 55.780 48.340 ;
        RECT 50.440 48.030 55.780 48.090 ;
        RECT 50.440 47.720 56.630 48.030 ;
        RECT 70.740 47.770 71.140 51.020 ;
        RECT 83.770 50.870 84.580 51.140 ;
        RECT 85.390 50.870 86.200 51.680 ;
        RECT 87.280 51.410 87.550 51.680 ;
        RECT 87.280 51.140 87.820 51.410 ;
        RECT 87.010 50.870 87.820 51.140 ;
        RECT 83.770 49.790 87.820 50.870 ;
        RECT 84.040 49.250 87.550 49.790 ;
        RECT 84.580 48.980 87.010 49.250 ;
        RECT 84.580 48.710 86.740 48.980 ;
        RECT 51.270 47.420 57.480 47.720 ;
        RECT 51.270 47.360 58.340 47.420 ;
        RECT 52.100 47.140 58.340 47.360 ;
        RECT 70.530 47.370 71.140 47.770 ;
        RECT 52.100 47.010 59.200 47.140 ;
        RECT 52.940 46.860 59.200 47.010 ;
        RECT 52.940 46.670 60.060 46.860 ;
        RECT 53.780 46.600 60.060 46.670 ;
        RECT 53.780 46.350 60.920 46.600 ;
        RECT 53.780 46.340 61.790 46.350 ;
        RECT 54.630 46.110 61.790 46.340 ;
        RECT 54.630 46.030 62.660 46.110 ;
        RECT 55.480 45.880 62.660 46.030 ;
        RECT 55.480 45.720 63.540 45.880 ;
        RECT 56.340 45.660 63.540 45.720 ;
        RECT 56.340 45.450 64.420 45.660 ;
        RECT 56.340 45.420 65.300 45.450 ;
        RECT 57.200 45.250 65.300 45.420 ;
        RECT 57.200 45.140 66.180 45.250 ;
        RECT 58.060 45.070 66.180 45.140 ;
        RECT 58.060 44.890 67.070 45.070 ;
        RECT 58.060 44.860 67.950 44.890 ;
        RECT 58.920 44.730 67.950 44.860 ;
        RECT 58.920 44.600 68.840 44.730 ;
        RECT 59.790 44.570 68.840 44.600 ;
        RECT 59.790 44.430 69.740 44.570 ;
        RECT 70.530 44.430 70.930 47.370 ;
        RECT 59.790 44.350 70.930 44.430 ;
        RECT 60.660 44.300 70.930 44.350 ;
        RECT 60.660 44.180 71.520 44.300 ;
        RECT 88.570 44.180 88.970 49.680 ;
        RECT 106.010 48.670 106.410 53.660 ;
        RECT 116.470 53.410 120.780 53.810 ;
        RECT 115.700 53.310 120.780 53.410 ;
        RECT 115.700 52.960 120.010 53.310 ;
        RECT 114.910 52.820 120.010 52.960 ;
        RECT 114.910 52.520 119.250 52.820 ;
        RECT 114.120 52.340 119.250 52.520 ;
        RECT 114.120 52.090 118.470 52.340 ;
        RECT 113.330 51.870 118.470 52.090 ;
        RECT 113.330 51.670 117.700 51.870 ;
        RECT 112.520 51.410 117.700 51.670 ;
        RECT 112.520 51.260 116.910 51.410 ;
        RECT 111.720 50.960 116.910 51.260 ;
        RECT 111.720 50.860 116.120 50.960 ;
        RECT 110.910 50.520 116.120 50.860 ;
        RECT 110.910 50.470 115.330 50.520 ;
        RECT 110.090 50.090 115.330 50.470 ;
        RECT 109.270 49.720 114.520 50.090 ;
        RECT 108.440 49.670 114.520 49.720 ;
        RECT 108.440 49.360 113.720 49.670 ;
        RECT 107.610 49.260 113.720 49.360 ;
        RECT 107.610 49.010 112.910 49.260 ;
        RECT 106.780 48.860 112.910 49.010 ;
        RECT 106.780 48.670 112.090 48.860 ;
        RECT 105.940 48.470 112.090 48.670 ;
        RECT 105.940 48.340 111.270 48.470 ;
        RECT 105.100 48.090 111.270 48.340 ;
        RECT 105.100 48.030 110.440 48.090 ;
        RECT 104.250 47.720 110.440 48.030 ;
        RECT 103.400 47.420 109.610 47.720 ;
        RECT 102.540 47.360 109.610 47.420 ;
        RECT 102.540 47.140 108.780 47.360 ;
        RECT 101.680 47.010 108.780 47.140 ;
        RECT 101.680 46.860 107.940 47.010 ;
        RECT 100.820 46.670 107.940 46.860 ;
        RECT 100.820 46.600 107.100 46.670 ;
        RECT 99.960 46.350 107.100 46.600 ;
        RECT 99.090 46.340 107.100 46.350 ;
        RECT 99.090 46.110 106.250 46.340 ;
        RECT 98.220 46.030 106.250 46.110 ;
        RECT 98.220 45.880 105.400 46.030 ;
        RECT 97.340 45.720 105.400 45.880 ;
        RECT 97.340 45.660 104.540 45.720 ;
        RECT 96.460 45.450 104.540 45.660 ;
        RECT 95.580 45.420 104.540 45.450 ;
        RECT 95.580 45.250 103.680 45.420 ;
        RECT 94.700 45.140 103.680 45.250 ;
        RECT 94.700 45.070 102.820 45.140 ;
        RECT 93.810 44.890 102.820 45.070 ;
        RECT 92.930 44.860 102.820 44.890 ;
        RECT 92.930 44.730 101.960 44.860 ;
        RECT 92.040 44.600 101.960 44.730 ;
        RECT 92.040 44.570 101.090 44.600 ;
        RECT 91.140 44.430 101.090 44.570 ;
        RECT 90.250 44.350 101.090 44.430 ;
        RECT 90.250 44.300 100.220 44.350 ;
        RECT 89.360 44.180 100.220 44.300 ;
        RECT 60.660 44.110 72.420 44.180 ;
        RECT 61.540 44.070 72.420 44.110 ;
        RECT 88.460 44.110 100.220 44.180 ;
        RECT 88.460 44.070 99.340 44.110 ;
        RECT 61.540 43.980 73.320 44.070 ;
        RECT 87.560 43.980 99.340 44.070 ;
        RECT 61.540 43.890 74.220 43.980 ;
        RECT 86.660 43.890 99.340 43.980 ;
        RECT 61.540 43.880 75.120 43.890 ;
        RECT 62.420 43.820 75.120 43.880 ;
        RECT 85.760 43.880 99.340 43.890 ;
        RECT 85.760 43.820 98.460 43.880 ;
        RECT 62.420 43.760 76.020 43.820 ;
        RECT 84.860 43.760 98.460 43.820 ;
        RECT 62.420 43.710 76.920 43.760 ;
        RECT 83.960 43.710 98.460 43.760 ;
        RECT 62.420 43.670 77.830 43.710 ;
        RECT 83.050 43.670 98.460 43.710 ;
        RECT 62.420 43.660 78.730 43.670 ;
        RECT 63.300 43.640 78.730 43.660 ;
        RECT 82.150 43.660 98.460 43.670 ;
        RECT 82.150 43.640 97.580 43.660 ;
        RECT 63.300 43.620 79.640 43.640 ;
        RECT 81.240 43.620 97.580 43.640 ;
        RECT 63.300 43.450 97.580 43.620 ;
        RECT 64.180 43.250 96.700 43.450 ;
        RECT 65.070 43.070 95.810 43.250 ;
        RECT 65.950 42.890 94.930 43.070 ;
        RECT 66.840 42.730 94.040 42.890 ;
        RECT 67.740 42.570 93.140 42.730 ;
        RECT 68.630 42.430 92.250 42.570 ;
        RECT 69.520 42.300 91.360 42.430 ;
        RECT 70.420 42.180 90.460 42.300 ;
        RECT 71.320 42.070 89.560 42.180 ;
        RECT 72.220 41.980 88.660 42.070 ;
        RECT 73.120 41.890 87.760 41.980 ;
        RECT 74.020 41.820 86.860 41.890 ;
        RECT 74.920 41.760 85.960 41.820 ;
        RECT 75.830 41.710 85.050 41.760 ;
        RECT 76.730 41.670 84.150 41.710 ;
        RECT 77.640 41.640 83.240 41.670 ;
        RECT 78.540 41.620 82.340 41.640 ;
        RECT 79.440 41.610 81.430 41.620 ;
      LAYER met3 ;
        RECT 85.810 223.665 86.230 224.265 ;
        RECT 88.570 223.665 88.990 224.265 ;
        RECT 91.330 223.665 91.750 224.265 ;
        RECT 91.720 221.360 92.300 221.370 ;
        RECT 90.300 219.400 90.800 220.000 ;
        RECT 61.410 218.030 62.100 218.730 ;
        RECT 91.560 217.050 92.560 221.360 ;
        RECT 85.360 216.050 92.560 217.050 ;
      LAYER met3 ;
        RECT 34.060 149.220 40.260 162.320 ;
        RECT 48.050 160.370 54.250 173.470 ;
        RECT 64.690 166.900 70.890 180.000 ;
        RECT 82.520 168.240 88.720 181.340 ;
      LAYER met3 ;
        RECT 90.270 174.670 90.890 175.140 ;
      LAYER met3 ;
        RECT 99.960 164.260 106.160 177.360 ;
        RECT 115.440 155.310 121.640 168.410 ;
      LAYER met3 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 68.170 149.600 91.570 152.200 ;
      LAYER met3 ;
        RECT 23.990 134.440 30.190 147.540 ;
      LAYER met3 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 60.370 134.000 99.370 144.400 ;
      LAYER met3 ;
        RECT 127.610 142.200 133.810 155.300 ;
      LAYER met3 ;
        RECT 60.370 131.400 68.170 134.000 ;
      LAYER met3 ;
        RECT 18.870 117.350 25.070 130.450 ;
      LAYER met3 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
      LAYER met3 ;
        RECT 135.520 126.090 141.720 139.190 ;
      LAYER met3 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 0.530 114.410 2.770 114.870 ;
        RECT 7.470 114.410 9.070 114.435 ;
        RECT 0.530 112.910 9.070 114.410 ;
        RECT 30.710 114.305 31.810 115.555 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 0.530 112.330 2.770 112.910 ;
        RECT 7.470 112.885 9.070 112.910 ;
      LAYER met3 ;
        RECT 18.720 99.470 24.920 112.570 ;
      LAYER met3 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
      LAYER met3 ;
        RECT 138.040 108.410 144.240 121.510 ;
      LAYER met3 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
      LAYER met3 ;
        RECT 24.140 82.380 30.340 95.480 ;
      LAYER met3 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
      LAYER met3 ;
        RECT 135.520 90.730 141.720 103.830 ;
      LAYER met3 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
      LAYER met3 ;
        RECT 34.210 67.400 40.410 80.500 ;
      LAYER met3 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
      LAYER met3 ;
        RECT 127.760 74.620 133.960 87.720 ;
        RECT 48.190 56.250 54.390 69.350 ;
        RECT 64.840 49.720 71.040 62.820 ;
        RECT 82.670 48.380 88.870 61.480 ;
        RECT 100.110 52.360 106.310 65.460 ;
        RECT 115.590 61.310 121.790 74.410 ;
      LAYER met4 ;
        RECT 30.670 223.050 30.970 224.760 ;
        RECT 33.430 223.050 33.730 224.760 ;
        RECT 36.190 223.050 36.490 224.760 ;
        RECT 38.950 223.050 39.250 224.760 ;
        RECT 41.710 223.050 42.010 224.760 ;
        RECT 44.470 223.050 44.770 224.760 ;
        RECT 47.230 223.050 47.530 224.760 ;
        RECT 49.990 223.050 50.290 224.760 ;
        RECT 52.750 223.050 53.050 224.760 ;
        RECT 55.510 223.050 55.810 224.760 ;
        RECT 58.270 223.050 58.570 224.760 ;
        RECT 61.030 223.050 61.330 224.760 ;
        RECT 63.790 223.050 64.090 224.760 ;
        RECT 66.550 223.050 66.850 224.760 ;
        RECT 69.310 223.050 69.610 224.760 ;
        RECT 72.070 223.050 72.370 224.760 ;
        RECT 74.830 223.050 75.130 224.760 ;
        RECT 77.590 223.050 77.890 224.760 ;
        RECT 80.350 223.050 80.650 224.760 ;
        RECT 83.110 223.050 83.410 224.760 ;
        RECT 85.870 224.095 86.170 224.760 ;
        RECT 88.630 224.095 88.930 224.760 ;
        RECT 91.390 224.095 91.690 224.760 ;
        RECT 85.855 223.685 86.185 224.095 ;
        RECT 88.615 223.685 88.945 224.095 ;
        RECT 91.375 223.685 91.705 224.095 ;
        RECT 1.000 222.050 83.410 223.050 ;
        RECT 94.150 222.110 94.450 224.760 ;
        RECT 1.000 220.760 2.500 222.050 ;
        RECT 60.490 218.650 61.490 222.050 ;
        RECT 90.410 221.810 94.450 222.110 ;
        RECT 90.410 220.000 90.710 221.810 ;
        RECT 90.300 219.400 90.800 220.000 ;
        RECT 60.490 218.140 62.030 218.650 ;
        RECT 61.490 218.110 62.030 218.140 ;
        RECT 85.405 217.050 86.415 217.055 ;
        RECT 5.500 216.050 86.415 217.050 ;
        RECT 85.405 216.045 86.415 216.050 ;
        RECT 90.410 175.145 90.710 219.400 ;
        RECT 90.315 174.665 90.845 175.145 ;
        RECT 90.410 174.640 90.710 174.665 ;
        RECT 70.770 152.200 91.570 154.800 ;
        RECT 68.170 149.600 91.570 152.200 ;
        RECT 62.970 144.400 96.770 149.600 ;
        RECT 60.370 134.000 99.370 144.400 ;
        RECT 60.370 131.400 68.170 134.000 ;
        RECT 60.370 128.800 65.570 131.400 ;
        RECT 62.970 126.200 65.570 128.800 ;
        RECT 75.970 126.200 83.770 134.000 ;
        RECT 91.570 131.400 99.370 134.000 ;
        RECT 94.170 128.800 99.370 131.400 ;
        RECT 94.170 126.200 96.770 128.800 ;
        RECT 62.970 123.600 68.170 126.200 ;
        RECT 73.370 123.600 86.370 126.200 ;
        RECT 91.570 123.600 96.770 126.200 ;
        RECT 62.970 121.000 78.570 123.600 ;
        RECT 81.170 121.000 94.170 123.600 ;
        RECT 68.170 118.400 75.970 121.000 ;
        RECT 83.770 118.400 94.170 121.000 ;
        RECT 0.575 112.325 1.000 114.875 ;
        RECT 2.500 112.325 2.725 114.875 ;
        RECT 5.500 114.110 31.920 115.610 ;
        RECT 70.770 113.200 88.970 118.400 ;
        RECT 55.170 110.600 62.970 113.200 ;
        RECT 70.770 110.600 73.370 113.200 ;
        RECT 75.970 110.600 78.570 113.200 ;
        RECT 81.170 110.600 83.770 113.200 ;
        RECT 86.370 110.600 88.970 113.200 ;
        RECT 96.770 110.600 104.570 113.200 ;
        RECT 52.570 105.400 65.570 110.600 ;
        RECT 94.170 105.400 107.170 110.600 ;
        RECT 55.170 102.800 70.770 105.400 ;
        RECT 88.970 102.800 104.570 105.400 ;
        RECT 62.970 100.200 73.370 102.800 ;
        RECT 86.370 100.200 96.770 102.800 ;
        RECT 68.170 97.600 78.570 100.200 ;
        RECT 81.170 97.600 91.570 100.200 ;
        RECT 73.370 92.400 86.370 97.600 ;
        RECT 68.170 89.800 78.570 92.400 ;
        RECT 81.170 89.800 91.570 92.400 ;
        RECT 55.170 87.200 73.370 89.800 ;
        RECT 86.370 87.200 107.170 89.800 ;
        RECT 52.570 84.600 68.170 87.200 ;
        RECT 91.570 84.600 107.170 87.200 ;
        RECT 52.570 82.000 62.970 84.600 ;
        RECT 96.770 82.000 107.170 84.600 ;
        RECT 52.570 79.400 60.370 82.000 ;
        RECT 99.370 79.400 107.170 82.000 ;
        RECT 55.170 76.800 57.770 79.400 ;
        RECT 101.970 76.800 104.570 79.400 ;
  END
END tt_um_oscillating_bones
END LIBRARY

