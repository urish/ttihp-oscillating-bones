* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] ua[0] ua[1] ua[2] ua[3] ua[4] ua[5] ua[6] ua[7] VAPWR
+ VDPWR VGND
X0 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VAPWR.t15 VAPWR.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X1 VGND.t35 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_5.A VGND.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X2 VDPWR.t61 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_10715_43723# VDPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X3 a_10297_43723# a_10168_43997# a_9876_43697# VGND.t53 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X4 a_10544_44089# a_10297_43723# VDPWR.t45 VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X5 uo_out[0].t1 ua[0].t2 VGND.t47 VGND.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X6 a_10368_43697# a_10161_43697# a_10544_44089# VDPWR.t51 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X7 VGND.t65 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X8 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VAPWR.t33 VAPWR.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X9 VGND.t51 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X10 ua[0].t1 skullfet_3v3_buffer.A VAPWR.t25 VAPWR.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X11 a_13468_43697# a_13740_43697# VGND.t75 VGND.t74 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X12 VDPWR.t31 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12647_43723# VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X13 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VAPWR.t35 VAPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X14 a_14232_43697# a_14032_43997# a_14381_43723# VGND.t103 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X15 VGND.t7 a_11441_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t6 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X16 VAPWR.t5 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VAPWR.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X17 a_12093_43697# uo_out[1].t2 VDPWR.t37 VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X18 a_12051_44089# a_11536_43697# VDPWR.t13 VDPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X19 VAPWR.t7 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VAPWR.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X20 VGND.t117 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X21 VGND.t5 a_13468_43697# uo_out[1].t1 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X22 VDPWR.t73 a_9509_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VDPWR.t72 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X23 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VGND.t25 VGND.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X24 ring_0/skullfet_inverter_9.A skullfet_3v3_buffer.A VAPWR.t23 VAPWR.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X25 a_13960_43723# a_13468_43697# VGND.t3 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X26 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t113 VGND.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X27 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t37 VGND.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X28 VGND.t43 a_9604_43697# uo_out[3].t1 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X29 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t115 VGND.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X30 VAPWR.t13 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VAPWR.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X31 VGND.t77 a_14232_43697# a_14161_43723# VGND.t76 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X32 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VAPWR.t19 VAPWR.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X33 VGND.t87 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X34 VGND.t107 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X35 a_12647_43723# a_12100_43997# a_12300_43697# VDPWR.t57 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X36 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t73 VGND.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X37 a_13468_43697# a_13740_43697# VDPWR.t53 VDPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X38 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VAPWR.t31 VAPWR.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X39 a_11441_43697# a_11536_43697# VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X40 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t21 VGND.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X41 VDPWR.t50 a_10161_43697# a_10168_43997# VDPWR.t49 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X42 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_5.A VAPWR.t27 VAPWR.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X43 a_14025_43697# uo_out[0].t2 VGND.t27 VGND.t26 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X44 a_14232_43697# a_14025_43697# a_14408_44089# VDPWR.t65 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X45 a_14161_43723# a_14025_43697# a_13740_43697# VDPWR.t64 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X46 VDPWR.t5 a_13468_43697# uo_out[1].t0 VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X47 VDPWR.t17 a_12093_43697# a_12100_43997# VDPWR.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X48 VDPWR.t29 a_9604_43697# uo_out[3].t0 VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X49 VGND.t95 a_14025_43697# a_14032_43997# VGND.t94 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X50 a_9509_43697# a_9604_43697# VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X51 VGND.t109 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X52 a_10119_44089# a_9604_43697# VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X53 a_10161_43697# uo_out[2].t2 VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X54 a_13740_43697# a_14032_43997# a_13983_44089# VDPWR.t71 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X55 VAPWR.t21 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VAPWR.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X56 VGND.t97 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X57 a_12028_43723# a_11536_43697# VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X58 skullfet_3v3_buffer.A ring_0/skullfet_inverter_7.A VAPWR.t17 VAPWR.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X59 a_10517_43723# a_10297_43723# VGND.t63 VGND.t62 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X60 VAPWR.t41 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VAPWR.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X61 VGND.t83 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_6.A VGND.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X62 a_9604_43697# a_9876_43697# VGND.t101 VGND.t100 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X63 VGND.t89 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_14579_43723# VGND.t88 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X64 a_12093_43697# uo_out[1].t3 VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X65 VAPWR.t3 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VAPWR.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X66 a_12449_43723# a_12229_43723# VGND.t61 VGND.t60 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X67 VGND.t13 a_11536_43697# uo_out[2].t1 VGND.t12 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X68 VGND.t111 a_9509_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t110 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X69 VGND.t105 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t104 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X70 VGND.t99 a_12300_43697# a_12229_43723# VGND.t98 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X71 a_10715_43723# a_10168_43997# a_10368_43697# VDPWR.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X72 a_9604_43697# a_9876_43697# VDPWR.t69 VDPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X73 a_11536_43697# a_11808_43697# VDPWR.t39 VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X74 a_13373_43697# a_13468_43697# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X75 a_14408_44089# a_14161_43723# VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X76 VGND.t55 ring_0/skullfet_inverter_7.A skullfet_3v3_buffer.A VGND.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X77 VGND.t71 a_10161_43697# a_10168_43997# VGND.t70 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X78 a_10096_43723# a_9604_43697# VGND.t41 VGND.t40 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X79 VDPWR.t35 ua[0].t3 uo_out[0].t0 VDPWR.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X80 VDPWR.t9 a_11536_43697# uo_out[2].t0 VDPWR.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X81 VDPWR.t41 a_13373_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X82 a_14579_43723# a_14025_43697# a_14232_43697# VGND.t93 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X83 a_14161_43723# a_14032_43997# a_13740_43697# VGND.t102 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X84 VDPWR.t59 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_14579_43723# VDPWR.t58 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X85 VGND.t19 a_12093_43697# a_12100_43997# VGND.t18 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X86 a_10368_43697# a_10168_43997# a_10517_43723# VGND.t52 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X87 a_11808_43697# a_12100_43997# a_12051_44089# VDPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X88 VAPWR.t11 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VAPWR.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X89 a_10161_43697# uo_out[2].t3 VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X90 VAPWR.t39 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VAPWR.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=5.3775 pd=12.07 as=7.5825 ps=29.53 w=4.5 l=0.5
X91 a_11536_43697# a_11808_43697# VGND.t57 VGND.t56 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X92 a_12300_43697# a_12100_43997# a_12449_43723# VGND.t85 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X93 a_11808_43697# a_12093_43697# a_12028_43723# VGND.t17 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X94 VGND.t67 a_10368_43697# a_10297_43723# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X95 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VAPWR.t1 VAPWR.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X96 a_13373_43697# a_13468_43697# VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X97 a_13740_43697# a_14025_43697# a_13960_43723# VGND.t92 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X98 VDPWR.t55 a_14232_43697# a_14161_43723# VDPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X99 a_10297_43723# a_10161_43697# a_9876_43697# VDPWR.t48 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X100 VGND.t81 skullfet_3v3_buffer.A ua[0].t0 VGND.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X101 a_12229_43723# a_12100_43997# a_11808_43697# VGND.t84 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X102 a_11441_43697# a_11536_43697# VGND.t11 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X103 a_12476_44089# a_12229_43723# VDPWR.t43 VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X104 a_10715_43723# a_10161_43697# a_10368_43697# VGND.t69 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X105 a_12229_43723# a_12093_43697# a_11808_43697# VDPWR.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X106 a_12300_43697# a_12093_43697# a_12476_44089# VDPWR.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X107 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VAPWR.t29 VAPWR.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X108 VDPWR.t7 a_11441_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X109 VGND.t9 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X110 VGND.t79 skullfet_3v3_buffer.A ring_0/skullfet_inverter_9.A VGND.t78 sky130_fd_pr__nfet_g5v0d10v5 ad=5.1075 pd=11.95 as=7.8525 ps=29.65 w=4.5 l=0.5
X111 VGND.t59 a_13373_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X112 a_12647_43723# a_12093_43697# a_12300_43697# VGND.t16 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X113 a_9509_43697# a_9604_43697# VGND.t39 VGND.t38 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X114 VGND.t91 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_10715_43723# VGND.t90 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X115 a_9876_43697# a_10168_43997# a_10119_44089# VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X116 ring_0/skullfet_inverter_5.A ring_0/skullfet_inverter_4.A VAPWR.t9 VAPWR.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X117 a_14381_43723# a_14161_43723# VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X118 VGND.t45 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_12647_43723# VGND.t44 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X119 a_14579_43723# a_14032_43997# a_14232_43697# VDPWR.t70 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X120 a_9876_43697# a_10161_43697# a_10096_43723# VGND.t68 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X121 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VGND.t23 VGND.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X122 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VAPWR.t37 VAPWR.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X123 VDPWR.t47 a_10368_43697# a_10297_43723# VDPWR.t46 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X124 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VAPWR.t43 VAPWR.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=7.5825 pd=29.53 as=5.3775 ps=12.07 w=4.5 l=0.5
X125 a_14025_43697# uo_out[0].t3 VDPWR.t19 VDPWR.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X126 a_13983_44089# a_13468_43697# VDPWR.t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X127 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t49 VGND.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=7.8525 pd=29.65 as=5.1075 ps=11.95 w=4.5 l=0.5
X128 VDPWR.t67 a_12300_43697# a_12229_43723# VDPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X129 VDPWR.t63 a_14025_43697# a_14032_43997# VDPWR.t62 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
R0 VAPWR.n66 VAPWR.t25 738.801
R1 VAPWR.n52 VAPWR.t21 738.799
R2 VAPWR.n54 VAPWR.t19 738.799
R3 VAPWR.n38 VAPWR.t5 738.799
R4 VAPWR.n34 VAPWR.t7 738.799
R5 VAPWR.n6 VAPWR.t31 738.799
R6 VAPWR.n41 VAPWR.t41 738.799
R7 VAPWR.n44 VAPWR.t11 738.799
R8 VAPWR.n47 VAPWR.t39 738.799
R9 VAPWR.n4 VAPWR.t3 738.799
R10 VAPWR.n2 VAPWR.t13 738.799
R11 VAPWR.n60 VAPWR.t37 738.799
R12 VAPWR.n57 VAPWR.t29 738.799
R13 VAPWR.n32 VAPWR.t1 738.799
R14 VAPWR.n7 VAPWR.t35 738.799
R15 VAPWR.n11 VAPWR.t27 738.799
R16 VAPWR.n22 VAPWR.t15 738.799
R17 VAPWR.n19 VAPWR.t17 738.799
R18 VAPWR.n16 VAPWR.t23 738.799
R19 VAPWR.n13 VAPWR.t43 738.799
R20 VAPWR.n9 VAPWR.t9 738.799
R21 VAPWR.n27 VAPWR.t33 738.799
R22 VAPWR.n60 VAPWR.t36 707.519
R23 VAPWR.n57 VAPWR.t28 707.519
R24 VAPWR.n52 VAPWR.t20 707.519
R25 VAPWR.n54 VAPWR.t18 707.519
R26 VAPWR.n38 VAPWR.t4 707.519
R27 VAPWR.n34 VAPWR.t6 707.519
R28 VAPWR.n32 VAPWR.t0 707.519
R29 VAPWR.n6 VAPWR.t30 707.519
R30 VAPWR.n7 VAPWR.t34 707.519
R31 VAPWR.n11 VAPWR.t26 707.519
R32 VAPWR.n22 VAPWR.t14 707.519
R33 VAPWR.n19 VAPWR.t16 707.519
R34 VAPWR.n16 VAPWR.t22 707.519
R35 VAPWR.n13 VAPWR.t42 707.519
R36 VAPWR.n9 VAPWR.t8 707.519
R37 VAPWR.n27 VAPWR.t32 707.519
R38 VAPWR.n41 VAPWR.t40 707.519
R39 VAPWR.n44 VAPWR.t10 707.519
R40 VAPWR.n47 VAPWR.t38 707.519
R41 VAPWR.n4 VAPWR.t2 707.519
R42 VAPWR.n2 VAPWR.t12 707.519
R43 VAPWR.n66 VAPWR.t24 707.519
R44 VAPWR.n67 VAPWR 13.899
R45 VAPWR.n61 VAPWR.n60 13.3797
R46 VAPWR.n58 VAPWR.n57 13.3797
R47 VAPWR.n33 VAPWR.n32 13.3797
R48 VAPWR.n8 VAPWR.n7 13.3797
R49 VAPWR.n12 VAPWR.n11 13.3797
R50 VAPWR.n23 VAPWR.n22 13.3797
R51 VAPWR.n20 VAPWR.n19 13.3797
R52 VAPWR.n17 VAPWR.n16 13.3797
R53 VAPWR.n14 VAPWR.n13 13.3797
R54 VAPWR.n10 VAPWR.n9 13.3797
R55 VAPWR.n28 VAPWR.n27 13.3797
R56 VAPWR.n53 VAPWR.n52 13.3223
R57 VAPWR VAPWR.n54 13.3223
R58 VAPWR.n39 VAPWR.n38 13.3223
R59 VAPWR.n35 VAPWR.n34 13.3223
R60 VAPWR VAPWR.n6 13.3223
R61 VAPWR.n42 VAPWR.n41 13.3223
R62 VAPWR.n45 VAPWR.n44 13.3223
R63 VAPWR.n48 VAPWR.n47 13.3223
R64 VAPWR.n5 VAPWR.n4 13.3223
R65 VAPWR.n3 VAPWR.n2 13.3223
R66 VAPWR VAPWR.n66 13.3223
R67 VAPWR.n59 VAPWR.n58 9.70762
R68 VAPWR.n18 VAPWR.n15 9.45042
R69 VAPWR.n31 VAPWR 8.52916
R70 VAPWR.n62 VAPWR.n61 7.92611
R71 VAPWR.n40 VAPWR.n37 7.71912
R72 VAPWR.n15 VAPWR.n14 7.71771
R73 VAPWR.n31 VAPWR.n30 7.41572
R74 VAPWR.n55 VAPWR 7.13154
R75 VAPWR.n40 VAPWR.n39 7.11663
R76 VAPWR.n18 VAPWR.n17 7.10884
R77 VAPWR.n43 VAPWR.n42 6.89753
R78 VAPWR.n21 VAPWR.n20 6.54898
R79 VAPWR.n49 VAPWR.n46 6.23852
R80 VAPWR.n30 VAPWR.n8 6.19396
R81 VAPWR.n46 VAPWR.n45 6.10554
R82 VAPWR.n29 VAPWR.n28 6.01845
R83 VAPWR.n36 VAPWR.n35 5.92055
R84 VAPWR.n49 VAPWR.n48 5.84717
R85 VAPWR.n24 VAPWR.n23 5.78073
R86 VAPWR.n26 VAPWR.n10 5.73072
R87 VAPWR.n50 VAPWR.n5 5.60146
R88 VAPWR.n51 VAPWR.n3 5.59565
R89 VAPWR.n25 VAPWR.n12 5.50466
R90 VAPWR.n55 VAPWR.n53 4.89777
R91 VAPWR.n36 VAPWR.n33 4.86074
R92 VAPWR.n46 VAPWR.n43 4.01511
R93 VAPWR.n67 VAPWR 3.49636
R94 VAPWR.n69 VAPWR 3.44936
R95 VAPWR.n37 VAPWR.n36 2.91269
R96 VAPWR.n59 VAPWR.n56 2.82184
R97 VAPWR.n1 VAPWR.n0 1.63622
R98 VAPWR.n24 VAPWR.n21 1.36014
R99 VAPWR.n30 VAPWR.n29 1.34127
R100 VAPWR.n56 VAPWR.n51 1.32921
R101 VAPWR.n56 VAPWR.n55 1.313
R102 VAPWR.n63 VAPWR.n0 1.29727
R103 VAPWR.n29 VAPWR.n26 1.10191
R104 VAPWR.n51 VAPWR.n50 0.940035
R105 VAPWR.n62 VAPWR.n59 0.85748
R106 VAPWR.n37 VAPWR.n31 0.767594
R107 VAPWR.n68 VAPWR.n65 0.616014
R108 VAPWR.n25 VAPWR.n24 0.52495
R109 VAPWR.n43 VAPWR.n40 0.514977
R110 VAPWR.n15 VAPWR.n1 0.507476
R111 VAPWR.n26 VAPWR.n25 0.505442
R112 VAPWR.n21 VAPWR.n18 0.500622
R113 VAPWR.n50 VAPWR.n49 0.483622
R114 VAPWR.n65 VAPWR.n0 0.20333
R115 VAPWR VAPWR.n69 0.193138
R116 VAPWR.n61 VAPWR 0.057877
R117 VAPWR.n58 VAPWR 0.057877
R118 VAPWR.n33 VAPWR 0.057877
R119 VAPWR.n8 VAPWR 0.057877
R120 VAPWR.n12 VAPWR 0.057877
R121 VAPWR.n23 VAPWR 0.057877
R122 VAPWR.n20 VAPWR 0.057877
R123 VAPWR.n17 VAPWR 0.057877
R124 VAPWR.n14 VAPWR 0.057877
R125 VAPWR.n10 VAPWR 0.057877
R126 VAPWR.n28 VAPWR 0.057877
R127 VAPWR.n53 VAPWR 0.0496071
R128 VAPWR.n39 VAPWR 0.0496071
R129 VAPWR.n35 VAPWR 0.0496071
R130 VAPWR.n42 VAPWR 0.0496071
R131 VAPWR.n45 VAPWR 0.0496071
R132 VAPWR.n48 VAPWR 0.0496071
R133 VAPWR.n5 VAPWR 0.0496071
R134 VAPWR.n3 VAPWR 0.0496071
R135 VAPWR.n65 VAPWR.n64 0.0335189
R136 VAPWR.n64 VAPWR.n1 0.00474612
R137 VAPWR.n63 VAPWR.n62 0.00305102
R138 VAPWR.n64 VAPWR.n63 0.00285849
R139 VAPWR.n68 VAPWR.n67 0.0018126
R140 VAPWR.n69 VAPWR.n68 0.0018126
R141 VGND.n209 VGND.n194 101372
R142 VGND.n272 VGND.n158 97829.8
R143 VGND.n234 VGND.n183 63317.7
R144 VGND.n228 VGND.n217 49981.2
R145 VGND.n230 VGND.t108 48989.1
R146 VGND.n195 VGND.n182 48956.8
R147 VGND.n226 VGND.n159 34056.2
R148 VGND.n218 VGND.n118 31758
R149 VGND.n431 VGND.n52 31668.4
R150 VGND.n326 VGND.n325 31013.9
R151 VGND.n201 VGND.n196 31013.9
R152 VGND.n325 VGND.n324 30664.6
R153 VGND.n204 VGND.n196 30664.6
R154 VGND.n225 VGND.n224 30639.5
R155 VGND.n430 VGND.n53 29705.2
R156 VGND.n228 VGND.n184 26125.9
R157 VGND.n231 VGND.n230 24501.8
R158 VGND.n233 VGND.n184 22668.4
R159 VGND.n195 VGND.n194 20954.6
R160 VGND.n158 VGND.n53 20954.6
R161 VGND.n229 VGND.n193 18294.4
R162 VGND.n328 VGND.n52 16731.6
R163 VGND.n196 VGND.n195 13862.9
R164 VGND.n325 VGND.n53 13853.3
R165 VGND.n230 VGND.n184 10983.3
R166 VGND.n328 VGND.t98 10623.7
R167 VGND.t72 VGND.n234 8761.83
R168 VGND.n233 VGND.n232 8254.98
R169 VGND.n194 VGND.n183 8164.43
R170 VGND.n234 VGND.n233 8000.6
R171 VGND.n270 VGND.n160 7798.05
R172 VGND.n219 VGND.n218 7223.1
R173 VGND.n228 VGND.n183 6658.85
R174 VGND.n193 VGND.n187 6298.11
R175 VGND.n211 VGND.n160 6257.53
R176 VGND.n225 VGND.n158 6251.53
R177 VGND.n234 VGND.n182 5608.83
R178 VGND.n226 VGND.n225 4619.12
R179 VGND.n264 VGND.t8 4526.67
R180 VGND.n217 VGND.n210 4456.64
R181 VGND.n231 VGND.n185 4323.23
R182 VGND.n193 VGND.n192 4311.21
R183 VGND.n213 VGND.n211 3590.94
R184 VGND.n269 VGND.t8 3461.39
R185 VGND.n271 VGND.n159 3297.03
R186 VGND.n227 VGND.n160 3097.77
R187 VGND.n229 VGND.n228 3097.77
R188 VGND.n216 VGND.n214 3043.22
R189 VGND.n270 VGND.t106 2956.47
R190 VGND.n192 VGND.n191 2374.28
R191 VGND.n192 VGND.n189 2325.64
R192 VGND.n209 VGND.t114 2293.69
R193 VGND.n235 VGND.t72 2108.34
R194 VGND.n214 VGND.n160 2021.45
R195 VGND.n218 VGND.t110 1534.08
R196 VGND.n187 VGND.t116 1523.34
R197 VGND.t22 VGND.n216 1523.34
R198 VGND.n272 VGND.t104 1467.82
R199 VGND.n221 VGND.n219 1240.19
R200 VGND.t48 VGND.n182 1206.01
R201 VGND.n329 VGND.n76 1198.25
R202 VGND.n369 VGND.n368 1198.25
R203 VGND.n367 VGND.n63 1198.25
R204 VGND.n331 VGND.n330 1198.25
R205 VGND.n211 VGND.t8 1196.46
R206 VGND.t106 VGND.n159 1186.75
R207 VGND.n161 VGND.n159 921.593
R208 VGND.n208 VGND.n206 892.495
R209 VGND.t20 VGND.n198 842.21
R210 VGND.t18 VGND.t44 800.774
R211 VGND.t0 VGND.t4 797.881
R212 VGND.n273 VGND.t34 787.793
R213 VGND.n326 VGND.t50 779.42
R214 VGND.n118 VGND 684.976
R215 VGND.n272 VGND.n271 655.47
R216 VGND.n210 VGND.n209 634.295
R217 VGND.n224 VGND.n223 600.63
R218 VGND.n330 VGND.t58 596.322
R219 VGND.n221 VGND.n220 585
R220 VGND.n187 VGND.n186 585
R221 VGND.n189 VGND.n188 585
R222 VGND.n191 VGND.n190 585
R223 VGND.n323 VGND.n322 585
R224 VGND.n433 VGND.n432 585
R225 VGND.n295 VGND.n119 585
R226 VGND.n274 VGND.n273 585
R227 VGND.n200 VGND.n199 585
R228 VGND.n198 VGND.n197 585
R229 VGND.n203 VGND.n202 585
R230 VGND.n206 VGND.n205 585
R231 VGND.n208 VGND.n207 585
R232 VGND.n216 VGND.n215 585
R233 VGND.n213 VGND.n212 585
R234 VGND.n269 VGND.n268 585
R235 VGND.n223 VGND.n222 585
R236 VGND.n366 VGND.n365 585
R237 VGND.n428 VGND.n427 585
R238 VGND.n189 VGND.t108 574.539
R239 VGND.n324 VGND.t82 539.317
R240 VGND.t112 VGND.n201 533.332
R241 VGND.t36 VGND.n204 500.077
R242 VGND.t44 VGND.t16 477.058
R243 VGND.n431 VGND.n430 425.618
R244 VGND.n232 VGND.t64 424.175
R245 VGND.n327 VGND.n118 422.882
R246 VGND.t16 VGND.t85 421.685
R247 VGND.t85 VGND.t60 421.685
R248 VGND.n430 VGND.n429 405.947
R249 VGND.t58 VGND.t0 404.647
R250 VGND.n330 VGND.n329 391.868
R251 VGND.n329 VGND 391.868
R252 VGND.n201 VGND.n200 382.728
R253 VGND.t74 VGND.t2 381.911
R254 VGND.t56 VGND.t14 381.911
R255 VGND.n324 VGND.n119 377.945
R256 VGND.t94 VGND.t88 377.889
R257 VGND.t10 VGND.t12 377.889
R258 VGND.t70 VGND.t90 377.889
R259 VGND.t38 VGND.t42 377.889
R260 VGND.n191 VGND.t86 362.452
R261 VGND.n217 VGND.t22 360.884
R262 VGND.n204 VGND.n203 360.842
R263 VGND.t28 VGND.t18 357.793
R264 VGND.n273 VGND.n272 302.216
R265 VGND.n264 VGND.t9 282.13
R266 VGND.n161 VGND.t107 282.13
R267 VGND.n295 VGND.t35 282.13
R268 VGND.n433 VGND.t51 282.13
R269 VGND.n188 VGND.t109 282.13
R270 VGND.n220 VGND.t79 282.13
R271 VGND.n186 VGND.t117 282.13
R272 VGND.n190 VGND.t87 282.13
R273 VGND.n222 VGND.t55 282.13
R274 VGND.n322 VGND.t83 282.13
R275 VGND.n274 VGND.t105 282.13
R276 VGND.n365 VGND.t47 281.841
R277 VGND.n427 VGND.t81 281.841
R278 VGND.n235 VGND.t73 281.839
R279 VGND.n215 VGND.t23 281.839
R280 VGND.n212 VGND.t25 281.839
R281 VGND.n185 VGND.t65 281.839
R282 VGND.n268 VGND.t97 281.839
R283 VGND.n207 VGND.t115 281.839
R284 VGND.n205 VGND.t37 281.839
R285 VGND.n202 VGND.t113 281.839
R286 VGND.n197 VGND.t49 281.839
R287 VGND.n199 VGND.t21 281.839
R288 VGND.n368 VGND.t6 281.408
R289 VGND.n230 VGND.n229 264.286
R290 VGND.n107 VGND.t3 251
R291 VGND.n354 VGND.t15 251
R292 VGND.n392 VGND.t41 251
R293 VGND.n232 VGND.t86 245.631
R294 VGND.n94 VGND.t89 243.028
R295 VGND.n341 VGND.t45 243.028
R296 VGND.n379 VGND.t91 243.028
R297 VGND.t76 VGND.t32 239.196
R298 VGND.n429 VGND.t54 237.476
R299 VGND.t88 VGND.t93 225.126
R300 VGND.n432 VGND.t50 222.331
R301 VGND.n81 VGND.n80 218.506
R302 VGND.n68 VGND.n67 218.506
R303 VGND.n394 VGND.n393 218.506
R304 VGND.n224 VGND.t78 214.124
R305 VGND.t92 VGND.t102 213.065
R306 VGND.t17 VGND.t84 213.065
R307 VGND.t68 VGND.t53 213.065
R308 VGND.n228 VGND.n227 209.014
R309 VGND.t80 VGND.t40 205.025
R310 VGND.t102 VGND.t76 203.016
R311 VGND.n78 VGND.n77 200.201
R312 VGND.n65 VGND.n64 200.201
R313 VGND.n402 VGND.n401 200.201
R314 VGND.n90 VGND.n89 199.739
R315 VGND.n337 VGND.n336 199.739
R316 VGND.n375 VGND.n374 199.739
R317 VGND.n100 VGND.n85 199.53
R318 VGND.n347 VGND.n73 199.53
R319 VGND.n385 VGND.n60 199.53
R320 VGND.t32 VGND.t103 198.995
R321 VGND.t69 VGND.t52 198.995
R322 VGND.t52 VGND.t62 198.995
R323 VGND.n223 VGND.t54 196.702
R324 VGND.n429 VGND.t66 194.976
R325 VGND.t2 VGND.t92 190.956
R326 VGND.t14 VGND.t17 190.956
R327 VGND.t6 VGND.t10 190.956
R328 VGND.t40 VGND.t68 190.956
R329 VGND.t110 VGND.t38 190.956
R330 VGND.n368 VGND.n367 184.925
R331 VGND.n367 VGND.t46 182.916
R332 VGND.n366 VGND.t69 178.894
R333 VGND.n214 VGND.n210 178.196
R334 VGND.t100 VGND.t80 176.885
R335 VGND.t26 VGND.t94 168.845
R336 VGND.t4 VGND.t74 168.845
R337 VGND.t12 VGND.t56 168.845
R338 VGND.t30 VGND.t70 168.845
R339 VGND.t42 VGND.t100 168.845
R340 VGND.t78 VGND.n221 164.337
R341 VGND.t82 VGND.n323 162.868
R342 VGND.t34 VGND.n119 153.912
R343 VGND.n203 VGND.t112 153.888
R344 VGND.n200 VGND.t20 151.095
R345 VGND.n198 VGND.t48 151.095
R346 VGND.n206 VGND.t36 145.869
R347 VGND.t60 VGND.n328 136.303
R348 VGND VGND.t28 132.043
R349 VGND.n214 VGND.t24 130.082
R350 VGND.n270 VGND.t96 129.425
R351 VGND.n271 VGND.n270 127.109
R352 VGND.t66 VGND.n428 120.603
R353 VGND.n327 VGND.t93 118.594
R354 VGND.t24 VGND.n213 99.8351
R355 VGND.t96 VGND.n269 99.332
R356 VGND.n219 VGND.n193 93.5857
R357 VGND.n428 VGND.t53 82.4126
R358 VGND.t103 VGND.n327 80.4025
R359 VGND.n85 VGND.t77 74.8666
R360 VGND.n73 VGND.t99 74.8666
R361 VGND.n60 VGND.t67 74.8666
R362 VGND.n209 VGND.n208 73.7658
R363 VGND.t84 VGND.n52 72.3623
R364 VGND.n327 VGND.n326 66.8513
R365 VGND VGND.t26 62.3121
R366 VGND VGND.t30 62.3121
R367 VGND.t64 VGND.n231 54.4208
R368 VGND.n77 VGND.t1 54.2862
R369 VGND.n64 VGND.t11 54.2862
R370 VGND.n401 VGND.t39 54.2862
R371 VGND.n323 VGND.n118 53.7948
R372 VGND.t90 VGND.n366 46.2317
R373 VGND.n429 VGND.t62 44.2216
R374 VGND.n85 VGND.t33 40.0005
R375 VGND.n73 VGND.t61 40.0005
R376 VGND.n60 VGND.t63 40.0005
R377 VGND.n89 VGND.t27 38.5719
R378 VGND.n89 VGND.t95 38.5719
R379 VGND.n336 VGND.t29 38.5719
R380 VGND.n336 VGND.t19 38.5719
R381 VGND.n374 VGND.t31 38.5719
R382 VGND.n374 VGND.t71 38.5719
R383 VGND.n432 VGND.n431 34.9453
R384 VGND.n112 VGND.n111 34.6358
R385 VGND.n113 VGND.n112 34.6358
R386 VGND.n102 VGND.n101 34.6358
R387 VGND.n102 VGND.n83 34.6358
R388 VGND.n106 VGND.n83 34.6358
R389 VGND.n95 VGND.n87 34.6358
R390 VGND.n99 VGND.n87 34.6358
R391 VGND.n343 VGND.n342 34.6358
R392 VGND.n343 VGND.n72 34.6358
R393 VGND.n349 VGND.n348 34.6358
R394 VGND.n349 VGND.n70 34.6358
R395 VGND.n353 VGND.n70 34.6358
R396 VGND.n359 VGND.n358 34.6358
R397 VGND.n360 VGND.n359 34.6358
R398 VGND.n381 VGND.n380 34.6358
R399 VGND.n381 VGND.n59 34.6358
R400 VGND.n387 VGND.n386 34.6358
R401 VGND.n387 VGND.n57 34.6358
R402 VGND.n391 VGND.n57 34.6358
R403 VGND.n399 VGND.n55 34.6358
R404 VGND.n400 VGND.n399 34.6358
R405 VGND.n108 VGND.n81 32.7534
R406 VGND.n355 VGND.n68 32.7534
R407 VGND.n395 VGND.n394 32.7534
R408 VGND.n108 VGND.n107 31.2476
R409 VGND.n355 VGND.n354 31.2476
R410 VGND.n395 VGND.n392 31.2476
R411 VGND.n100 VGND.n99 30.8711
R412 VGND.n347 VGND.n72 30.8711
R413 VGND.n385 VGND.n59 30.8711
R414 VGND.n95 VGND.n94 27.4829
R415 VGND.n342 VGND.n341 27.4829
R416 VGND.n380 VGND.n379 27.4829
R417 VGND.n77 VGND.t59 25.9346
R418 VGND.n64 VGND.t7 25.9346
R419 VGND.n401 VGND.t111 25.9346
R420 VGND.n80 VGND.t75 24.9236
R421 VGND.n80 VGND.t5 24.9236
R422 VGND.n67 VGND.t57 24.9236
R423 VGND.n67 VGND.t13 24.9236
R424 VGND.n393 VGND.t101 24.9236
R425 VGND.n393 VGND.t43 24.9236
R426 VGND.n262 VGND.n261 23.8791
R427 VGND.n331 VGND.n117 23.7181
R428 VGND.n113 VGND.n78 23.7181
R429 VGND.n335 VGND.n76 23.7181
R430 VGND.n360 VGND.n65 23.7181
R431 VGND.n369 VGND.n364 23.7181
R432 VGND.n373 VGND.n63 23.7181
R433 VGND.n402 VGND.n400 23.7181
R434 VGND.n236 VGND.n1 23.1262
R435 VGND.n93 VGND.n90 22.9652
R436 VGND.n94 VGND.n93 22.9652
R437 VGND.n337 VGND.n75 22.9652
R438 VGND.n341 VGND.n75 22.9652
R439 VGND.n375 VGND.n62 22.9652
R440 VGND.n379 VGND.n62 22.9652
R441 VGND.n107 VGND.n106 22.2123
R442 VGND.n354 VGND.n353 22.2123
R443 VGND.n392 VGND.n391 22.2123
R444 VGND.n117 VGND.n78 21.4593
R445 VGND.n337 VGND.n335 21.4593
R446 VGND.n364 VGND.n65 21.4593
R447 VGND.n375 VGND.n373 21.4593
R448 VGND.n488 VGND.n487 20.8917
R449 VGND.n267 VGND.n163 19.445
R450 VGND.n227 VGND.n226 15.7795
R451 VGND.n265 VGND.n264 13.2958
R452 VGND.n162 VGND.n161 13.2958
R453 VGND.n296 VGND.n295 13.2958
R454 VGND.n434 VGND.n433 13.2958
R455 VGND.n188 VGND.n3 13.2958
R456 VGND.n220 VGND.n8 13.2958
R457 VGND.n186 VGND.n4 13.2958
R458 VGND.n190 VGND.n2 13.2958
R459 VGND.n222 VGND.n32 13.2958
R460 VGND.n322 VGND.n321 13.2958
R461 VGND.n275 VGND.n274 13.2958
R462 VGND.n365 VGND 13.2396
R463 VGND.n215 VGND 13.2396
R464 VGND.n212 VGND 13.2396
R465 VGND.n185 VGND 13.2396
R466 VGND.n268 VGND 13.2396
R467 VGND.n207 VGND 13.2396
R468 VGND.n205 VGND 13.2396
R469 VGND.n197 VGND 13.2396
R470 VGND.n199 VGND 13.2396
R471 VGND.n202 VGND 13.2396
R472 VGND VGND.n235 13.2396
R473 VGND.n427 VGND 13.2396
R474 VGND.n331 VGND.n76 12.8005
R475 VGND.n369 VGND.n63 12.8005
R476 VGND.n263 VGND.n262 11.3685
R477 VGND.n101 VGND.n100 10.5417
R478 VGND.n348 VGND.n347 10.5417
R479 VGND.n386 VGND.n385 10.5417
R480 VGND.n400 VGND.n54 9.3005
R481 VGND.n399 VGND.n398 9.3005
R482 VGND.n397 VGND.n55 9.3005
R483 VGND.n396 VGND.n395 9.3005
R484 VGND.n392 VGND.n56 9.3005
R485 VGND.n391 VGND.n390 9.3005
R486 VGND.n389 VGND.n57 9.3005
R487 VGND.n388 VGND.n387 9.3005
R488 VGND.n386 VGND.n58 9.3005
R489 VGND.n385 VGND.n384 9.3005
R490 VGND.n383 VGND.n59 9.3005
R491 VGND.n382 VGND.n381 9.3005
R492 VGND.n380 VGND.n61 9.3005
R493 VGND.n379 VGND.n378 9.3005
R494 VGND.n377 VGND.n62 9.3005
R495 VGND.n376 VGND.n375 9.3005
R496 VGND.n373 VGND.n372 9.3005
R497 VGND.n371 VGND.n63 9.3005
R498 VGND.n93 VGND.n92 9.3005
R499 VGND.n94 VGND.n88 9.3005
R500 VGND.n96 VGND.n95 9.3005
R501 VGND.n97 VGND.n87 9.3005
R502 VGND.n99 VGND.n98 9.3005
R503 VGND.n100 VGND.n86 9.3005
R504 VGND.n101 VGND.n84 9.3005
R505 VGND.n103 VGND.n102 9.3005
R506 VGND.n104 VGND.n83 9.3005
R507 VGND.n106 VGND.n105 9.3005
R508 VGND.n107 VGND.n82 9.3005
R509 VGND.n109 VGND.n108 9.3005
R510 VGND.n111 VGND.n110 9.3005
R511 VGND.n112 VGND.n79 9.3005
R512 VGND.n114 VGND.n113 9.3005
R513 VGND.n115 VGND.n78 9.3005
R514 VGND.n117 VGND.n116 9.3005
R515 VGND.n333 VGND.n76 9.3005
R516 VGND.n335 VGND.n334 9.3005
R517 VGND.n338 VGND.n337 9.3005
R518 VGND.n339 VGND.n75 9.3005
R519 VGND.n341 VGND.n340 9.3005
R520 VGND.n342 VGND.n74 9.3005
R521 VGND.n344 VGND.n343 9.3005
R522 VGND.n345 VGND.n72 9.3005
R523 VGND.n347 VGND.n346 9.3005
R524 VGND.n348 VGND.n71 9.3005
R525 VGND.n350 VGND.n349 9.3005
R526 VGND.n351 VGND.n70 9.3005
R527 VGND.n353 VGND.n352 9.3005
R528 VGND.n354 VGND.n69 9.3005
R529 VGND.n356 VGND.n355 9.3005
R530 VGND.n358 VGND.n357 9.3005
R531 VGND.n359 VGND.n66 9.3005
R532 VGND.n361 VGND.n360 9.3005
R533 VGND.n362 VGND.n65 9.3005
R534 VGND.n364 VGND.n363 9.3005
R535 VGND.n370 VGND.n369 9.3005
R536 VGND.n332 VGND.n331 9.3005
R537 VGND VGND.n1 9.06372
R538 VGND.n266 VGND.n265 7.80496
R539 VGND.n163 VGND.n162 7.42221
R540 VGND.n91 VGND.n90 7.12576
R541 VGND.n403 VGND.n402 7.12063
R542 VGND.n425 VGND.n424 7.0515
R543 VGND.n489 VGND.n3 6.96
R544 VGND.n236 VGND 6.82321
R545 VGND.n490 VGND.n2 6.32363
R546 VGND.n276 VGND.n275 6.24462
R547 VGND VGND.n181 6.10287
R548 VGND VGND.n267 5.99098
R549 VGND.n262 VGND 5.98182
R550 VGND.n488 VGND.n4 5.94997
R551 VGND.n482 VGND.n8 5.91022
R552 VGND.n261 VGND 5.81859
R553 VGND.n321 VGND.n320 5.80858
R554 VGND.n297 VGND.n296 5.70662
R555 VGND.n257 VGND 5.69376
R556 VGND.n260 VGND 5.57954
R557 VGND.n259 VGND 5.53239
R558 VGND.n263 VGND 5.49935
R559 VGND.n458 VGND.n32 5.39911
R560 VGND.n424 VGND.n0 5.35255
R561 VGND.n319 VGND.n121 5.04217
R562 VGND.n435 VGND.n434 5.00883
R563 VGND.n426 VGND 4.99008
R564 VGND VGND.n426 4.97064
R565 VGND.n425 VGND 4.76873
R566 VGND.n0 VGND 3.44325
R567 VGND.n493 VGND 3.36335
R568 VGND.n319 VGND.n318 3.29217
R569 VGND.n163 VGND.n157 3.10947
R570 VGND VGND.n493 2.3855
R571 VGND.t46 VGND 2.01055
R572 VGND.n111 VGND.n81 1.88285
R573 VGND.n358 VGND.n68 1.88285
R574 VGND.n394 VGND.n55 1.88285
R575 VGND.n469 VGND.n468 1.5618
R576 VGND.n426 VGND.n425 1.44737
R577 VGND.n266 VGND.n263 1.28628
R578 VGND.n435 VGND.n50 1.2755
R579 VGND.n320 VGND.n120 0.979021
R580 VGND.n237 VGND.n236 0.96878
R581 VGND.n490 VGND.n489 0.964749
R582 VGND.n267 VGND.n266 0.93288
R583 VGND.n489 VGND.n488 0.903134
R584 VGND.n260 VGND.n259 0.844578
R585 VGND.n470 VGND.n469 0.777168
R586 VGND.n492 VGND.n491 0.726602
R587 VGND.n261 VGND.n260 0.707232
R588 VGND.n320 VGND.n319 0.6755
R589 VGND.n436 VGND.n435 0.638
R590 VGND.n259 VGND.n258 0.577069
R591 VGND.n315 VGND.n120 0.574766
R592 VGND.n491 VGND.n1 0.561048
R593 VGND.n471 VGND.n470 0.533644
R594 VGND.n315 VGND.n314 0.469554
R595 VGND.n314 VGND.n313 0.431514
R596 VGND.n318 VGND.n51 0.425271
R597 VGND.n472 VGND.n471 0.420347
R598 VGND.n404 uo_out[4] 0.4094
R599 VGND.n405 uo_out[5] 0.4094
R600 VGND.n406 uo_out[6] 0.4094
R601 VGND.n407 uo_out[7] 0.4094
R602 VGND.n408 uio_out[0] 0.4094
R603 VGND.n409 uio_out[1] 0.4094
R604 VGND.n410 uio_out[2] 0.4094
R605 VGND.n411 uio_out[3] 0.4094
R606 uio_out[5] VGND.n421 0.4094
R607 uio_out[6] VGND.n420 0.4094
R608 uio_out[7] VGND.n419 0.4094
R609 uio_oe[0] VGND.n418 0.4094
R610 uio_oe[1] VGND.n417 0.4094
R611 uio_oe[2] VGND.n416 0.4094
R612 uio_oe[3] VGND.n415 0.4094
R613 uio_oe[4] VGND.n414 0.4094
R614 uio_oe[5] VGND.n413 0.4094
R615 uio_oe[6] VGND.n412 0.4094
R616 VGND.n473 VGND.n472 0.36938
R617 VGND.n313 VGND.n312 0.355217
R618 VGND.n474 VGND.n473 0.332442
R619 VGND.n312 VGND.n311 0.314827
R620 VGND.n258 VGND.n164 0.307815
R621 VGND.n475 VGND.n474 0.293921
R622 VGND.n423 VGND.n422 0.284067
R623 VGND.n311 VGND.n310 0.283145
R624 VGND.n424 VGND.n423 0.2684
R625 VGND.n476 VGND.n475 0.262603
R626 VGND.n310 VGND.n309 0.257575
R627 VGND.n477 VGND.n476 0.242676
R628 VGND.n309 VGND.n308 0.242107
R629 VGND.n478 VGND.n477 0.227688
R630 VGND.n308 VGND.n307 0.224203
R631 VGND.n297 VGND.n294 0.21925
R632 VGND.n479 VGND.n478 0.214493
R633 VGND.n307 VGND.n306 0.209128
R634 VGND.n238 VGND.n237 0.207265
R635 VGND.n479 VGND.n11 0.207112
R636 VGND.n478 VGND.n12 0.205418
R637 VGND.n477 VGND.n13 0.203752
R638 VGND.n254 VGND.n164 0.202174
R639 VGND.n480 VGND.n479 0.201991
R640 VGND.n476 VGND.n14 0.2005
R641 VGND.n475 VGND.n15 0.198913
R642 VGND.n474 VGND.n16 0.19735
R643 VGND.n306 VGND.n305 0.196195
R644 VGND.n473 VGND.n17 0.195812
R645 VGND.n481 VGND.n480 0.194723
R646 VGND.n472 VGND.n18 0.194298
R647 VGND.n483 VGND.n482 0.193682
R648 VGND.n471 VGND.n19 0.19134
R649 VGND.n254 VGND.n253 0.190823
R650 VGND.n470 VGND.n20 0.189894
R651 VGND.n305 VGND.n304 0.189066
R652 VGND.n469 VGND.n21 0.18847
R653 VGND.n487 VGND.n5 0.188059
R654 VGND.n253 VGND.n252 0.184664
R655 VGND.n486 VGND.n485 0.181056
R656 VGND.n252 VGND.n251 0.180457
R657 VGND.n304 VGND.n303 0.179109
R658 VGND.n303 VGND.n302 0.178762
R659 VGND.n251 VGND.n250 0.167949
R660 VGND.n302 VGND.n301 0.166149
R661 VGND.n276 VGND.n157 0.165057
R662 VGND.n249 VGND.n248 0.164532
R663 VGND.n250 VGND.n249 0.164276
R664 VGND.n300 VGND.n299 0.159573
R665 VGND.n301 VGND.n300 0.159247
R666 VGND.n441 VGND.n440 0.159247
R667 VGND.n460 VGND.n459 0.156646
R668 VGND.n442 VGND.n441 0.156448
R669 VGND.n248 VGND.n247 0.155102
R670 VGND.n316 VGND.n315 0.154588
R671 VGND.n480 VGND.n10 0.153861
R672 VGND.n314 VGND.n122 0.153802
R673 VGND.n299 VGND.n298 0.153257
R674 VGND.n247 VGND.n246 0.153062
R675 VGND.n313 VGND.n123 0.153016
R676 VGND VGND.n403 0.152603
R677 VGND.n440 VGND.n50 0.152527
R678 VGND.n311 VGND.n125 0.152399
R679 VGND.n436 VGND.n51 0.152332
R680 VGND.n312 VGND.n124 0.15223
R681 VGND.n444 VGND.n443 0.151068
R682 VGND.n309 VGND.n127 0.150816
R683 VGND.n246 VGND.n245 0.150802
R684 VGND.n310 VGND.n126 0.150657
R685 VGND.n443 VGND.n442 0.15035
R686 VGND.n307 VGND.n129 0.150182
R687 VGND.n239 VGND.n179 0.150148
R688 VGND.n308 VGND.n128 0.150025
R689 VGND.n256 VGND.n164 0.149538
R690 VGND.n306 VGND.n130 0.149385
R691 VGND.n253 VGND.n165 0.148887
R692 VGND.n255 VGND.n254 0.148737
R693 VGND.n305 VGND.n131 0.148589
R694 VGND.n403 VGND.n54 0.148519
R695 VGND.n252 VGND.n166 0.148081
R696 VGND.n303 VGND.n133 0.147936
R697 VGND.n304 VGND.n132 0.147793
R698 VGND.n249 VGND.n169 0.147559
R699 VGND.n317 VGND.n121 0.147513
R700 VGND.n250 VGND.n168 0.147416
R701 VGND.n301 VGND.n135 0.147274
R702 VGND.n440 VGND.n439 0.147274
R703 VGND.n251 VGND.n167 0.147274
R704 VGND.n302 VGND.n134 0.147135
R705 VGND.n438 VGND.n437 0.147135
R706 VGND.n246 VGND.n172 0.147023
R707 VGND.n467 VGND.n23 0.146955
R708 VGND.n248 VGND.n170 0.146742
R709 VGND.n300 VGND.n136 0.146468
R710 VGND.n441 VGND.n49 0.146468
R711 VGND.n245 VGND.n173 0.146195
R712 VGND.n245 VGND.n244 0.146195
R713 VGND.n294 VGND.n293 0.146191
R714 VGND.n445 VGND.n444 0.146191
R715 VGND.n294 VGND.n139 0.145925
R716 VGND.n444 VGND.n46 0.145925
R717 VGND.n247 VGND.n171 0.145925
R718 VGND.n298 VGND.n138 0.145792
R719 VGND.n443 VGND.n47 0.145792
R720 VGND.n241 VGND.n177 0.14577
R721 VGND.n240 VGND.n178 0.14577
R722 VGND.n299 VGND.n137 0.145661
R723 VGND.n442 VGND.n48 0.145661
R724 VGND.n242 VGND.n176 0.145634
R725 VGND.n465 VGND.n25 0.145573
R726 VGND.n243 VGND.n175 0.1455
R727 VGND.n464 VGND.n26 0.145428
R728 VGND.n291 VGND.n142 0.145368
R729 VGND.n447 VGND.n43 0.145368
R730 VGND.n244 VGND.n174 0.145368
R731 VGND.n463 VGND.n27 0.145284
R732 VGND.n293 VGND.n140 0.145108
R733 VGND.n445 VGND.n45 0.145108
R734 VGND.n279 VGND.n154 0.144866
R735 VGND.n287 VGND.n146 0.144795
R736 VGND.n451 VGND.n39 0.144795
R737 VGND.n244 VGND.n243 0.144667
R738 VGND.n466 VGND.n24 0.144661
R739 VGND.n290 VGND.n143 0.14454
R740 VGND.n448 VGND.n42 0.14454
R741 VGND.n282 VGND.n151 0.144466
R742 VGND.n283 VGND.n150 0.144336
R743 VGND.n455 VGND.n35 0.144336
R744 VGND.n292 VGND.n141 0.144291
R745 VGND.n446 VGND.n44 0.144291
R746 VGND.n462 VGND.n28 0.14425
R747 VGND.n461 VGND.n29 0.144117
R748 VGND.n277 VGND.n156 0.144117
R749 VGND.n285 VGND.n148 0.144081
R750 VGND.n286 VGND.n147 0.144081
R751 VGND.n453 VGND.n37 0.144081
R752 VGND.n452 VGND.n38 0.144081
R753 VGND.n278 VGND.n155 0.143986
R754 VGND.n460 VGND.n30 0.143986
R755 VGND.n288 VGND.n145 0.143833
R756 VGND.n450 VGND.n40 0.143833
R757 VGND.n280 VGND.n153 0.143729
R758 VGND.n289 VGND.n144 0.143712
R759 VGND.n449 VGND.n41 0.143712
R760 VGND.n281 VGND.n152 0.143603
R761 VGND.n92 VGND.n91 0.143396
R762 VGND.n284 VGND.n149 0.143357
R763 VGND.n454 VGND.n36 0.143357
R764 VGND.n243 VGND.n242 0.143343
R765 VGND.n292 VGND.n291 0.142608
R766 VGND.n447 VGND.n446 0.142608
R767 VGND.n242 VGND.n241 0.142204
R768 VGND.n293 VGND.n292 0.14174
R769 VGND.n446 VGND.n445 0.14174
R770 VGND.n238 VGND.n180 0.141228
R771 VGND.n240 VGND.n239 0.140944
R772 VGND.n241 VGND.n240 0.14022
R773 VGND.n239 VGND.n238 0.139918
R774 VGND.n291 VGND.n290 0.138984
R775 VGND.n448 VGND.n447 0.138984
R776 VGND.n288 VGND.n287 0.137868
R777 VGND.n290 VGND.n289 0.137764
R778 VGND.n289 VGND.n288 0.13669
R779 VGND.n451 VGND.n450 0.135675
R780 VGND.n449 VGND.n448 0.135449
R781 VGND.n467 VGND.n466 0.134751
R782 VGND.n450 VGND.n449 0.134458
R783 VGND.n286 VGND.n285 0.134444
R784 VGND.n284 VGND.n283 0.13348
R785 VGND.n466 VGND.n465 0.133147
R786 VGND.n453 VGND.n452 0.132395
R787 VGND.n287 VGND.n286 0.132323
R788 VGND.n452 VGND.n451 0.132323
R789 VGND.n282 VGND.n281 0.131889
R790 VGND.n279 VGND.n278 0.131852
R791 VGND.n463 VGND.n462 0.13184
R792 VGND.n278 VGND.n277 0.131755
R793 VGND.n465 VGND.n464 0.131611
R794 VGND.n280 VGND.n279 0.131576
R795 VGND.n455 VGND.n454 0.131557
R796 VGND.n285 VGND.n284 0.131307
R797 VGND.n464 VGND.n463 0.131251
R798 VGND.n283 VGND.n282 0.130509
R799 VGND.n456 VGND.n455 0.130509
R800 VGND.n462 VGND.n461 0.130342
R801 VGND.n281 VGND.n280 0.130162
R802 VGND.n461 VGND.n460 0.13011
R803 VGND.n457 VGND.n456 0.130051
R804 VGND.n454 VGND.n453 0.129353
R805 VGND.n423 uio_out[4] 0.125833
R806 VGND.n23 VGND.n22 0.124567
R807 VGND.n92 VGND.n88 0.120292
R808 VGND.n96 VGND.n88 0.120292
R809 VGND.n97 VGND.n96 0.120292
R810 VGND.n98 VGND.n97 0.120292
R811 VGND.n98 VGND.n86 0.120292
R812 VGND.n86 VGND.n84 0.120292
R813 VGND.n103 VGND.n84 0.120292
R814 VGND.n104 VGND.n103 0.120292
R815 VGND.n105 VGND.n104 0.120292
R816 VGND.n105 VGND.n82 0.120292
R817 VGND.n109 VGND.n82 0.120292
R818 VGND.n110 VGND.n109 0.120292
R819 VGND.n110 VGND.n79 0.120292
R820 VGND.n114 VGND.n79 0.120292
R821 VGND.n115 VGND.n114 0.120292
R822 VGND.n116 VGND.n115 0.120292
R823 VGND.n339 VGND.n338 0.120292
R824 VGND.n340 VGND.n339 0.120292
R825 VGND.n340 VGND.n74 0.120292
R826 VGND.n344 VGND.n74 0.120292
R827 VGND.n345 VGND.n344 0.120292
R828 VGND.n346 VGND.n345 0.120292
R829 VGND.n346 VGND.n71 0.120292
R830 VGND.n350 VGND.n71 0.120292
R831 VGND.n351 VGND.n350 0.120292
R832 VGND.n352 VGND.n351 0.120292
R833 VGND.n352 VGND.n69 0.120292
R834 VGND.n356 VGND.n69 0.120292
R835 VGND.n357 VGND.n356 0.120292
R836 VGND.n357 VGND.n66 0.120292
R837 VGND.n361 VGND.n66 0.120292
R838 VGND.n362 VGND.n361 0.120292
R839 VGND.n363 VGND.n362 0.120292
R840 VGND.n377 VGND.n376 0.120292
R841 VGND.n378 VGND.n377 0.120292
R842 VGND.n378 VGND.n61 0.120292
R843 VGND.n382 VGND.n61 0.120292
R844 VGND.n383 VGND.n382 0.120292
R845 VGND.n384 VGND.n383 0.120292
R846 VGND.n384 VGND.n58 0.120292
R847 VGND.n388 VGND.n58 0.120292
R848 VGND.n389 VGND.n388 0.120292
R849 VGND.n390 VGND.n389 0.120292
R850 VGND.n390 VGND.n56 0.120292
R851 VGND.n396 VGND.n56 0.120292
R852 VGND.n397 VGND.n396 0.120292
R853 VGND.n398 VGND.n397 0.120292
R854 VGND.n398 VGND.n54 0.120292
R855 VGND.n456 VGND.n34 0.115155
R856 VGND.n437 VGND.n436 0.110794
R857 VGND.n12 VGND.n11 0.110004
R858 VGND.n459 VGND.n31 0.109215
R859 VGND.n13 VGND.n12 0.108082
R860 VGND.n14 VGND.n13 0.105175
R861 VGND.n157 VGND.n156 0.105059
R862 VGND.n11 VGND.n10 0.104833
R863 VGND.n468 VGND.n22 0.104045
R864 VGND.n15 VGND.n14 0.1015
R865 VGND.n16 VGND.n15 0.0997064
R866 VGND.n338 VGND 0.0981562
R867 VGND.n376 VGND 0.0981562
R868 VGND.n17 VGND.n16 0.097941
R869 VGND.n18 VGND.n17 0.0952266
R870 VGND.n33 VGND.n31 0.0946901
R871 VGND.n19 VGND.n18 0.0925543
R872 VGND.n486 VGND.n6 0.0910095
R873 VGND.n20 VGND.n19 0.0892405
R874 VGND.n21 VGND.n20 0.0876212
R875 VGND.n483 VGND.n6 0.0867209
R876 VGND.n7 VGND.n5 0.0867069
R877 VGND.n22 VGND.n21 0.0860263
R878 VGND.n468 VGND.n467 0.0819653
R879 VGND.n24 VGND.n23 0.0807239
R880 VGND.n458 VGND.n457 0.0803467
R881 VGND.n485 VGND.n5 0.0798478
R882 VGND.n484 VGND.n483 0.0787609
R883 VGND.n482 VGND.n7 0.0782778
R884 VGND.n481 VGND.n9 0.0776277
R885 VGND.n25 VGND.n24 0.0771423
R886 VGND.n26 VGND.n25 0.0762299
R887 VGND.n91 VGND 0.0758148
R888 VGND.n27 VGND.n26 0.0738696
R889 VGND.n9 VGND.n6 0.0721983
R890 VGND.n318 VGND.n317 0.0721201
R891 VGND.n487 VGND.n486 0.0720511
R892 VGND.n28 VGND.n27 0.0715432
R893 VGND.n29 VGND.n28 0.0701429
R894 VGND.n459 VGND.n458 0.0683371
R895 VGND.n30 VGND.n29 0.0678759
R896 VGND.n156 VGND.n155 0.0678759
R897 VGND.n35 VGND.n34 0.0675348
R898 VGND.n155 VGND.n154 0.0656408
R899 VGND.n31 VGND.n30 0.0656408
R900 VGND.n154 VGND.n153 0.0638803
R901 VGND.n153 VGND.n152 0.0621319
R902 VGND.n116 VGND 0.0603958
R903 VGND.n332 VGND 0.0603958
R904 VGND.n333 VGND 0.0603958
R905 VGND.n334 VGND 0.0603958
R906 VGND.n363 VGND 0.0603958
R907 VGND.n370 VGND 0.0603958
R908 VGND.n371 VGND 0.0603958
R909 VGND.n372 VGND 0.0603958
R910 VGND.n152 VGND.n151 0.0591207
R911 VGND.n10 VGND.n9 0.0590106
R912 VGND.n151 VGND.n150 0.0582586
R913 VGND.n265 VGND 0.05675
R914 VGND.n162 VGND 0.05675
R915 VGND.n296 VGND 0.05675
R916 VGND.n434 VGND 0.05675
R917 VGND.n3 VGND 0.05675
R918 VGND.n8 VGND 0.05675
R919 VGND.n4 VGND 0.05675
R920 VGND.n2 VGND 0.05675
R921 VGND.n32 VGND 0.05675
R922 VGND.n321 VGND 0.05675
R923 VGND.n275 VGND 0.05675
R924 VGND.n457 VGND.n33 0.0567284
R925 VGND.n150 VGND.n149 0.0561507
R926 VGND.n36 VGND.n35 0.0561507
R927 VGND.n149 VGND.n148 0.0549218
R928 VGND.n37 VGND.n36 0.0549218
R929 VGND.n180 VGND.n179 0.0533169
R930 VGND.n148 VGND.n147 0.0520203
R931 VGND.n38 VGND.n37 0.0520203
R932 VGND.n147 VGND.n146 0.0511757
R933 VGND.n39 VGND.n38 0.0511757
R934 VGND.n181 VGND.n180 0.0509967
R935 VGND.n179 VGND.n178 0.0486419
R936 VGND.n146 VGND.n145 0.0483188
R937 VGND.n40 VGND.n39 0.0483188
R938 VGND.n178 VGND.n177 0.0477973
R939 VGND.n404 uo_out[5] 0.0475
R940 VGND.n405 uo_out[6] 0.0475
R941 VGND.n406 uo_out[7] 0.0475
R942 VGND.n407 uio_out[0] 0.0475
R943 VGND.n408 uio_out[1] 0.0475
R944 VGND.n409 uio_out[2] 0.0475
R945 VGND.n410 uio_out[3] 0.0475
R946 VGND.n411 uio_out[4] 0.0475
R947 VGND.n422 uio_out[5] 0.0475
R948 VGND.n421 uio_out[6] 0.0475
R949 VGND.n420 uio_out[7] 0.0475
R950 VGND.n419 uio_oe[0] 0.0475
R951 VGND.n418 uio_oe[1] 0.0475
R952 VGND.n417 uio_oe[2] 0.0475
R953 VGND.n416 uio_oe[3] 0.0475
R954 VGND.n415 uio_oe[4] 0.0475
R955 VGND.n414 uio_oe[5] 0.0475
R956 VGND.n413 uio_oe[6] 0.0475
R957 VGND.n412 uio_oe[7] 0.0475
R958 VGND.n145 VGND.n144 0.0471667
R959 VGND.n41 VGND.n40 0.0471667
R960 VGND.n177 VGND.n176 0.045802
R961 VGND.n144 VGND.n143 0.045202
R962 VGND.n42 VGND.n41 0.045202
R963 VGND.n176 VGND.n175 0.0438333
R964 VGND.n143 VGND.n142 0.0435464
R965 VGND.n43 VGND.n42 0.0435464
R966 VGND.n142 VGND.n141 0.0418907
R967 VGND.n44 VGND.n43 0.0418907
R968 VGND.n175 VGND.n174 0.0418907
R969 VGND.n174 VGND.n173 0.0410629
R970 VGND.n484 VGND.n7 0.0407778
R971 VGND.n438 VGND.n51 0.0407077
R972 VGND.n141 VGND.n140 0.0405327
R973 VGND.n45 VGND.n44 0.0405327
R974 VGND.n173 VGND.n172 0.0385795
R975 VGND.n140 VGND.n139 0.0380817
R976 VGND.n46 VGND.n45 0.0380817
R977 VGND.n139 VGND.n138 0.0364477
R978 VGND.n47 VGND.n46 0.0364477
R979 VGND.n172 VGND.n171 0.0364477
R980 VGND.n171 VGND.n170 0.0356307
R981 VGND.n138 VGND.n137 0.0354026
R982 VGND.n48 VGND.n47 0.0354026
R983 VGND VGND.n332 0.0343542
R984 VGND VGND.n333 0.0343542
R985 VGND VGND.n370 0.0343542
R986 VGND VGND.n371 0.0343542
R987 VGND.n277 VGND.n276 0.0341879
R988 VGND.n170 VGND.n169 0.0331797
R989 VGND.n137 VGND.n136 0.0327581
R990 VGND.n49 VGND.n48 0.0327581
R991 VGND.n169 VGND.n168 0.0321558
R992 VGND.n136 VGND.n135 0.0319516
R993 VGND.n439 VGND.n49 0.0319516
R994 VGND.n34 VGND.n33 0.0307768
R995 VGND.n135 VGND.n134 0.0303387
R996 VGND.n439 VGND.n438 0.0303387
R997 VGND.n168 VGND.n167 0.0303387
R998 VGND.n482 VGND.n481 0.0297553
R999 VGND.n237 VGND.n181 0.0292963
R1000 VGND.n492 VGND.n0 0.0288333
R1001 VGND.n493 VGND.n492 0.0288333
R1002 VGND.n167 VGND.n166 0.0279194
R1003 VGND.n134 VGND.n133 0.0277436
R1004 VGND.n166 VGND.n165 0.0271129
R1005 VGND.n133 VGND.n132 0.0269423
R1006 VGND.n255 VGND.n165 0.0253397
R1007 VGND.n132 VGND.n131 0.0251815
R1008 uo_out[5] VGND.n404 0.024
R1009 uo_out[6] VGND.n405 0.024
R1010 uo_out[7] VGND.n406 0.024
R1011 uio_out[0] VGND.n407 0.024
R1012 uio_out[1] VGND.n408 0.024
R1013 uio_out[2] VGND.n409 0.024
R1014 uio_out[3] VGND.n410 0.024
R1015 uio_out[4] VGND.n411 0.024
R1016 VGND.n422 uio_out[5] 0.024
R1017 VGND.n421 uio_out[6] 0.024
R1018 VGND.n420 uio_out[7] 0.024
R1019 VGND.n419 uio_oe[0] 0.024
R1020 VGND.n418 uio_oe[1] 0.024
R1021 VGND.n417 uio_oe[2] 0.024
R1022 VGND.n416 uio_oe[3] 0.024
R1023 VGND.n415 uio_oe[4] 0.024
R1024 VGND.n414 uio_oe[5] 0.024
R1025 VGND.n413 uio_oe[6] 0.024
R1026 VGND.n412 uio_oe[7] 0.024
R1027 VGND.n256 VGND.n255 0.0237372
R1028 VGND.n131 VGND.n130 0.0235892
R1029 VGND.n334 VGND 0.0226354
R1030 VGND.n372 VGND 0.0226354
R1031 VGND.n130 VGND.n129 0.0219968
R1032 VGND.n257 VGND.n256 0.0219968
R1033 VGND.n129 VGND.n128 0.0204045
R1034 VGND.n128 VGND.n127 0.0186962
R1035 VGND.n298 VGND.n297 0.0175455
R1036 VGND.n127 VGND.n126 0.0171139
R1037 VGND.n126 VGND.n125 0.0154371
R1038 VGND.n437 VGND.n50 0.0141218
R1039 VGND.n125 VGND.n124 0.0139494
R1040 VGND.n485 VGND.n484 0.0135435
R1041 VGND.n124 VGND.n123 0.0122925
R1042 VGND.n123 VGND.n122 0.00993396
R1043 VGND.n258 VGND.n257 0.00918938
R1044 VGND.n316 VGND.n122 0.0091478
R1045 VGND.n317 VGND.n316 0.00757547
R1046 VGND.n121 VGND.n120 0.00689301
R1047 VGND.n491 VGND.n490 0.0011075
R1048 VDPWR.n1 VDPWR.t35 738.801
R1049 VDPWR.n1 VDPWR.t34 707.519
R1050 VDPWR.n84 VDPWR.t25 667.734
R1051 VDPWR.n52 VDPWR.t13 667.734
R1052 VDPWR.n124 VDPWR.t1 667.734
R1053 VDPWR.n99 VDPWR.t61 666.677
R1054 VDPWR.n38 VDPWR.t31 666.677
R1055 VDPWR.n4 VDPWR.t59 666.677
R1056 VDPWR.t52 VDPWR.t0 624.456
R1057 VDPWR.t12 VDPWR.t38 624.456
R1058 VDPWR.t24 VDPWR.t68 624.456
R1059 VDPWR.n102 VDPWR.n101 604.394
R1060 VDPWR.n33 VDPWR.n32 604.394
R1061 VDPWR.n142 VDPWR.n141 604.394
R1062 VDPWR.t58 VDPWR.t62 556.386
R1063 VDPWR.t2 VDPWR.t4 556.386
R1064 VDPWR.t16 VDPWR.t30 556.386
R1065 VDPWR.t8 VDPWR.t10 556.386
R1066 VDPWR.t49 VDPWR.t60 556.386
R1067 VDPWR.t28 VDPWR.t26 556.386
R1068 VDPWR.n17 VDPWR.t40 414.33
R1069 VDPWR.t6 VDPWR.n108 414.33
R1070 VDPWR.t54 VDPWR.t22 390.654
R1071 VDPWR.t42 VDPWR.t66 390.654
R1072 VDPWR.t44 VDPWR.t46 390.654
R1073 VDPWR.t0 VDPWR.t71 337.384
R1074 VDPWR.t56 VDPWR.t12 337.384
R1075 VDPWR.t32 VDPWR.t24 337.384
R1076 VDPWR.n82 VDPWR.n72 333.348
R1077 VDPWR.n54 VDPWR.n24 333.348
R1078 VDPWR.n122 VDPWR.n12 333.348
R1079 VDPWR.n68 VDPWR.n67 320.976
R1080 VDPWR.n45 VDPWR.n28 320.976
R1081 VDPWR.n9 VDPWR.n8 320.976
R1082 VDPWR.t22 VDPWR.t65 304.829
R1083 VDPWR.t14 VDPWR.t42 304.829
R1084 VDPWR.t51 VDPWR.t44 304.829
R1085 VDPWR.t40 VDPWR.t2 287.072
R1086 VDPWR.t10 VDPWR.t6 287.072
R1087 VDPWR.t26 VDPWR.t72 287.072
R1088 VDPWR.t65 VDPWR.t70 281.154
R1089 VDPWR.t64 VDPWR.t54 281.154
R1090 VDPWR.t57 VDPWR.t14 281.154
R1091 VDPWR.t66 VDPWR.t15 281.154
R1092 VDPWR.t33 VDPWR.t51 281.154
R1093 VDPWR.t46 VDPWR.t48 281.154
R1094 VDPWR.n109 VDPWR.n17 272.274
R1095 VDPWR.n109 VDPWR 272.274
R1096 VDPWR.n108 VDPWR.n107 272.274
R1097 VDPWR.n107 VDPWR 272.274
R1098 VDPWR.t70 VDPWR.t58 251.559
R1099 VDPWR.t30 VDPWR.t57 251.559
R1100 VDPWR.t60 VDPWR.t33 251.559
R1101 VDPWR.t62 VDPWR.t18 248.599
R1102 VDPWR.t71 VDPWR.t64 248.599
R1103 VDPWR.t4 VDPWR.t52 248.599
R1104 VDPWR.t36 VDPWR.t16 248.599
R1105 VDPWR.t15 VDPWR.t56 248.599
R1106 VDPWR.t38 VDPWR.t8 248.599
R1107 VDPWR.t20 VDPWR.t49 248.599
R1108 VDPWR.t48 VDPWR.t32 248.599
R1109 VDPWR.t68 VDPWR.t28 248.599
R1110 VDPWR.n76 VDPWR.n75 240.522
R1111 VDPWR.n60 VDPWR.n21 240.522
R1112 VDPWR.n116 VDPWR.n115 240.522
R1113 VDPWR.n107 VDPWR.n106 213.119
R1114 VDPWR.n108 VDPWR.n18 213.119
R1115 VDPWR.n110 VDPWR.n109 213.119
R1116 VDPWR.n17 VDPWR.n15 213.119
R1117 VDPWR.n67 VDPWR.t45 113.98
R1118 VDPWR.n28 VDPWR.t43 113.98
R1119 VDPWR.n8 VDPWR.t23 113.98
R1120 VDPWR.t18 VDPWR 91.745
R1121 VDPWR VDPWR.t36 91.745
R1122 VDPWR VDPWR.t20 91.745
R1123 VDPWR.n75 VDPWR.t27 61.9872
R1124 VDPWR.n21 VDPWR.t11 61.9872
R1125 VDPWR.n115 VDPWR.t3 61.9872
R1126 VDPWR.n101 VDPWR.t21 41.5552
R1127 VDPWR.n101 VDPWR.t50 41.5552
R1128 VDPWR.n32 VDPWR.t37 41.5552
R1129 VDPWR.n32 VDPWR.t17 41.5552
R1130 VDPWR.n141 VDPWR.t19 41.5552
R1131 VDPWR.n141 VDPWR.t63 41.5552
R1132 VDPWR.n67 VDPWR.t47 35.4605
R1133 VDPWR.n28 VDPWR.t67 35.4605
R1134 VDPWR.n8 VDPWR.t55 35.4605
R1135 VDPWR.n81 VDPWR.n73 34.6358
R1136 VDPWR.n77 VDPWR.n73 34.6358
R1137 VDPWR.n95 VDPWR.n65 34.6358
R1138 VDPWR.n95 VDPWR.n94 34.6358
R1139 VDPWR.n94 VDPWR.n93 34.6358
R1140 VDPWR.n90 VDPWR.n89 34.6358
R1141 VDPWR.n89 VDPWR.n88 34.6358
R1142 VDPWR.n88 VDPWR.n70 34.6358
R1143 VDPWR.n55 VDPWR.n22 34.6358
R1144 VDPWR.n59 VDPWR.n22 34.6358
R1145 VDPWR.n40 VDPWR.n39 34.6358
R1146 VDPWR.n40 VDPWR.n29 34.6358
R1147 VDPWR.n44 VDPWR.n29 34.6358
R1148 VDPWR.n47 VDPWR.n46 34.6358
R1149 VDPWR.n47 VDPWR.n26 34.6358
R1150 VDPWR.n51 VDPWR.n26 34.6358
R1151 VDPWR.n121 VDPWR.n13 34.6358
R1152 VDPWR.n117 VDPWR.n13 34.6358
R1153 VDPWR.n136 VDPWR.n135 34.6358
R1154 VDPWR.n135 VDPWR.n134 34.6358
R1155 VDPWR.n134 VDPWR.n6 34.6358
R1156 VDPWR.n130 VDPWR.n129 34.6358
R1157 VDPWR.n129 VDPWR.n128 34.6358
R1158 VDPWR.n128 VDPWR.n10 34.6358
R1159 VDPWR.n83 VDPWR.n82 32.0005
R1160 VDPWR.n54 VDPWR.n53 32.0005
R1161 VDPWR.n123 VDPWR.n122 32.0005
R1162 VDPWR.n143 VDPWR.n142 30.7593
R1163 VDPWR.n84 VDPWR.n83 30.4946
R1164 VDPWR.n53 VDPWR.n52 30.4946
R1165 VDPWR.n124 VDPWR.n123 30.4946
R1166 VDPWR.n75 VDPWR.t73 30.1692
R1167 VDPWR.n21 VDPWR.t7 30.1692
R1168 VDPWR.n115 VDPWR.t41 30.1692
R1169 VDPWR.n99 VDPWR.n65 27.4829
R1170 VDPWR.n61 VDPWR.n60 27.4829
R1171 VDPWR.n39 VDPWR.n38 27.4829
R1172 VDPWR.n116 VDPWR.n114 27.4829
R1173 VDPWR.n136 VDPWR.n4 27.4829
R1174 VDPWR.n72 VDPWR.t69 26.5955
R1175 VDPWR.n72 VDPWR.t29 26.5955
R1176 VDPWR.n24 VDPWR.t39 26.5955
R1177 VDPWR.n24 VDPWR.t9 26.5955
R1178 VDPWR.n12 VDPWR.t53 26.5955
R1179 VDPWR.n12 VDPWR.t5 26.5955
R1180 VDPWR.n77 VDPWR.n76 25.6005
R1181 VDPWR.n60 VDPWR.n59 25.6005
R1182 VDPWR.n117 VDPWR.n116 25.6005
R1183 VDPWR.n106 VDPWR.n19 23.7181
R1184 VDPWR.n61 VDPWR.n18 23.7181
R1185 VDPWR.n110 VDPWR.n16 23.7181
R1186 VDPWR.n114 VDPWR.n15 23.7181
R1187 VDPWR.n102 VDPWR.n100 22.9652
R1188 VDPWR.n37 VDPWR.n33 22.9652
R1189 VDPWR.n142 VDPWR.n140 22.9652
R1190 VDPWR.n100 VDPWR.n99 21.8358
R1191 VDPWR.n38 VDPWR.n37 21.8358
R1192 VDPWR.n140 VDPWR.n4 21.8358
R1193 VDPWR.n102 VDPWR.n19 21.4593
R1194 VDPWR.n33 VDPWR.n16 21.4593
R1195 VDPWR.n93 VDPWR.n68 18.4476
R1196 VDPWR.n45 VDPWR.n44 18.4476
R1197 VDPWR.n9 VDPWR.n6 18.4476
R1198 VDPWR.n90 VDPWR.n68 16.1887
R1199 VDPWR.n46 VDPWR.n45 16.1887
R1200 VDPWR.n130 VDPWR.n9 16.1887
R1201 VDPWR.n84 VDPWR.n70 15.0593
R1202 VDPWR.n52 VDPWR.n51 15.0593
R1203 VDPWR.n124 VDPWR.n10 15.0593
R1204 VDPWR.n2 VDPWR.n1 13.3223
R1205 VDPWR.n106 VDPWR.n18 12.8005
R1206 VDPWR.n110 VDPWR.n15 12.8005
R1207 VDPWR.n3 VDPWR 10.4834
R1208 VDPWR.n142 VDPWR.n0 9.3005
R1209 VDPWR.n140 VDPWR.n139 9.3005
R1210 VDPWR.n138 VDPWR.n4 9.3005
R1211 VDPWR.n137 VDPWR.n136 9.3005
R1212 VDPWR.n135 VDPWR.n5 9.3005
R1213 VDPWR.n134 VDPWR.n133 9.3005
R1214 VDPWR.n132 VDPWR.n6 9.3005
R1215 VDPWR.n131 VDPWR.n130 9.3005
R1216 VDPWR.n129 VDPWR.n7 9.3005
R1217 VDPWR.n128 VDPWR.n127 9.3005
R1218 VDPWR.n126 VDPWR.n10 9.3005
R1219 VDPWR.n125 VDPWR.n124 9.3005
R1220 VDPWR.n123 VDPWR.n11 9.3005
R1221 VDPWR.n121 VDPWR.n120 9.3005
R1222 VDPWR.n119 VDPWR.n13 9.3005
R1223 VDPWR.n118 VDPWR.n117 9.3005
R1224 VDPWR.n116 VDPWR.n14 9.3005
R1225 VDPWR.n114 VDPWR.n113 9.3005
R1226 VDPWR.n112 VDPWR.n15 9.3005
R1227 VDPWR.n111 VDPWR.n110 9.3005
R1228 VDPWR.n34 VDPWR.n16 9.3005
R1229 VDPWR.n35 VDPWR.n33 9.3005
R1230 VDPWR.n37 VDPWR.n36 9.3005
R1231 VDPWR.n38 VDPWR.n31 9.3005
R1232 VDPWR.n39 VDPWR.n30 9.3005
R1233 VDPWR.n41 VDPWR.n40 9.3005
R1234 VDPWR.n42 VDPWR.n29 9.3005
R1235 VDPWR.n44 VDPWR.n43 9.3005
R1236 VDPWR.n46 VDPWR.n27 9.3005
R1237 VDPWR.n48 VDPWR.n47 9.3005
R1238 VDPWR.n49 VDPWR.n26 9.3005
R1239 VDPWR.n51 VDPWR.n50 9.3005
R1240 VDPWR.n52 VDPWR.n25 9.3005
R1241 VDPWR.n53 VDPWR.n23 9.3005
R1242 VDPWR.n56 VDPWR.n55 9.3005
R1243 VDPWR.n57 VDPWR.n22 9.3005
R1244 VDPWR.n59 VDPWR.n58 9.3005
R1245 VDPWR.n60 VDPWR.n20 9.3005
R1246 VDPWR.n62 VDPWR.n61 9.3005
R1247 VDPWR.n63 VDPWR.n18 9.3005
R1248 VDPWR.n106 VDPWR.n105 9.3005
R1249 VDPWR.n104 VDPWR.n19 9.3005
R1250 VDPWR.n103 VDPWR.n102 9.3005
R1251 VDPWR.n100 VDPWR.n64 9.3005
R1252 VDPWR.n99 VDPWR.n98 9.3005
R1253 VDPWR.n97 VDPWR.n65 9.3005
R1254 VDPWR.n96 VDPWR.n95 9.3005
R1255 VDPWR.n94 VDPWR.n66 9.3005
R1256 VDPWR.n93 VDPWR.n92 9.3005
R1257 VDPWR.n91 VDPWR.n90 9.3005
R1258 VDPWR.n89 VDPWR.n69 9.3005
R1259 VDPWR.n88 VDPWR.n87 9.3005
R1260 VDPWR.n86 VDPWR.n70 9.3005
R1261 VDPWR.n85 VDPWR.n84 9.3005
R1262 VDPWR.n83 VDPWR.n71 9.3005
R1263 VDPWR.n81 VDPWR.n80 9.3005
R1264 VDPWR.n79 VDPWR.n73 9.3005
R1265 VDPWR.n78 VDPWR.n77 9.3005
R1266 VDPWR.n143 VDPWR.n3 8.8737
R1267 VDPWR.n76 VDPWR.n74 7.4049
R1268 VDPWR.n3 VDPWR.n2 6.49693
R1269 VDPWR.n82 VDPWR.n81 2.63579
R1270 VDPWR.n55 VDPWR.n54 2.63579
R1271 VDPWR.n122 VDPWR.n121 2.63579
R1272 VDPWR.n74 VDPWR 0.156264
R1273 VDPWR.n78 VDPWR.n74 0.144904
R1274 VDPWR.n139 VDPWR.n0 0.120292
R1275 VDPWR.n139 VDPWR.n138 0.120292
R1276 VDPWR.n138 VDPWR.n137 0.120292
R1277 VDPWR.n137 VDPWR.n5 0.120292
R1278 VDPWR.n133 VDPWR.n5 0.120292
R1279 VDPWR.n133 VDPWR.n132 0.120292
R1280 VDPWR.n132 VDPWR.n131 0.120292
R1281 VDPWR.n131 VDPWR.n7 0.120292
R1282 VDPWR.n127 VDPWR.n7 0.120292
R1283 VDPWR.n127 VDPWR.n126 0.120292
R1284 VDPWR.n126 VDPWR.n125 0.120292
R1285 VDPWR.n125 VDPWR.n11 0.120292
R1286 VDPWR.n120 VDPWR.n11 0.120292
R1287 VDPWR.n120 VDPWR.n119 0.120292
R1288 VDPWR.n119 VDPWR.n118 0.120292
R1289 VDPWR.n118 VDPWR.n14 0.120292
R1290 VDPWR.n113 VDPWR.n14 0.120292
R1291 VDPWR.n36 VDPWR.n35 0.120292
R1292 VDPWR.n36 VDPWR.n31 0.120292
R1293 VDPWR.n31 VDPWR.n30 0.120292
R1294 VDPWR.n41 VDPWR.n30 0.120292
R1295 VDPWR.n42 VDPWR.n41 0.120292
R1296 VDPWR.n43 VDPWR.n42 0.120292
R1297 VDPWR.n43 VDPWR.n27 0.120292
R1298 VDPWR.n48 VDPWR.n27 0.120292
R1299 VDPWR.n49 VDPWR.n48 0.120292
R1300 VDPWR.n50 VDPWR.n49 0.120292
R1301 VDPWR.n50 VDPWR.n25 0.120292
R1302 VDPWR.n25 VDPWR.n23 0.120292
R1303 VDPWR.n56 VDPWR.n23 0.120292
R1304 VDPWR.n57 VDPWR.n56 0.120292
R1305 VDPWR.n58 VDPWR.n57 0.120292
R1306 VDPWR.n58 VDPWR.n20 0.120292
R1307 VDPWR.n62 VDPWR.n20 0.120292
R1308 VDPWR.n103 VDPWR.n64 0.120292
R1309 VDPWR.n98 VDPWR.n64 0.120292
R1310 VDPWR.n98 VDPWR.n97 0.120292
R1311 VDPWR.n97 VDPWR.n96 0.120292
R1312 VDPWR.n96 VDPWR.n66 0.120292
R1313 VDPWR.n92 VDPWR.n66 0.120292
R1314 VDPWR.n92 VDPWR.n91 0.120292
R1315 VDPWR.n91 VDPWR.n69 0.120292
R1316 VDPWR.n87 VDPWR.n69 0.120292
R1317 VDPWR.n87 VDPWR.n86 0.120292
R1318 VDPWR.n86 VDPWR.n85 0.120292
R1319 VDPWR.n85 VDPWR.n71 0.120292
R1320 VDPWR.n80 VDPWR.n71 0.120292
R1321 VDPWR.n80 VDPWR.n79 0.120292
R1322 VDPWR.n79 VDPWR.n78 0.120292
R1323 VDPWR VDPWR.n0 0.0981562
R1324 VDPWR.n35 VDPWR 0.0981562
R1325 VDPWR VDPWR.n103 0.0981562
R1326 VDPWR.n113 VDPWR 0.0603958
R1327 VDPWR VDPWR.n112 0.0603958
R1328 VDPWR VDPWR.n111 0.0603958
R1329 VDPWR.n34 VDPWR 0.0603958
R1330 VDPWR VDPWR.n62 0.0603958
R1331 VDPWR.n63 VDPWR 0.0603958
R1332 VDPWR.n105 VDPWR 0.0603958
R1333 VDPWR VDPWR.n104 0.0603958
R1334 VDPWR.n2 VDPWR 0.0496071
R1335 VDPWR.n112 VDPWR 0.0382604
R1336 VDPWR.n111 VDPWR 0.0382604
R1337 VDPWR VDPWR.n63 0.0382604
R1338 VDPWR.n105 VDPWR 0.0382604
R1339 VDPWR VDPWR.n34 0.0226354
R1340 VDPWR.n104 VDPWR 0.0226354
R1341 VDPWR VDPWR.n143 0.0224072
R1342 ua[0] ua[0].t1 973.365
R1343 ua[0].n1 ua[0].t2 543.266
R1344 ua[0].n0 ua[0].t3 526.913
R1345 ua[0].n4 ua[0].t0 466.05
R1346 ua[0].n1 ua[0].n0 420.889
R1347 ua[0].n2 ua[0].n0 135.657
R1348 ua[0] ua[0].n1 117.829
R1349 ua[0].n3 ua[0] 48.4268
R1350 ua[0].n4 ua[0].n3 10.3749
R1351 ua[0].n2 ua[0] 10.2862
R1352 ua[0] ua[0].n4 10.0576
R1353 ua[0].n3 ua[0].n2 4.75847
R1354 uo_out[0].n0 uo_out[0].t0 983.422
R1355 uo_out[0] uo_out[0].t1 455.764
R1356 uo_out[0].n1 uo_out[0].t3 294.557
R1357 uo_out[0].n1 uo_out[0].t2 211.01
R1358 uo_out[0].n2 uo_out[0].n1 152
R1359 uo_out[0].n3 uo_out[0].n0 13.3264
R1360 uo_out[0].n3 uo_out[0].n2 13.1405
R1361 uo_out[0].n0 uo_out[0] 10.2862
R1362 uo_out[0].n4 uo_out[0] 8.14831
R1363 uo_out[0].n4 uo_out[0].n3 4.5005
R1364 uo_out[0].n2 uo_out[0] 2.01193
R1365 uo_out[0] uo_out[0].n4 0.0793043
R1366 uo_out[1].n2 uo_out[1].t0 313.104
R1367 uo_out[1].n0 uo_out[1].t2 294.557
R1368 uo_out[1].t1 uo_out[1].n2 265.769
R1369 uo_out[1] uo_out[1].t1 262.318
R1370 uo_out[1].n0 uo_out[1].t3 211.01
R1371 uo_out[1].n1 uo_out[1].n0 152
R1372 uo_out[1].n5 uo_out[1] 12.6752
R1373 uo_out[1].n4 uo_out[1].n1 11.6411
R1374 uo_out[1].n4 uo_out[1].n3 9.3005
R1375 uo_out[1].n3 uo_out[1] 7.17626
R1376 uo_out[1].n3 uo_out[1].n2 4.84898
R1377 uo_out[1].n5 uo_out[1].n4 4.5029
R1378 uo_out[1].n1 uo_out[1] 1.37896
R1379 uo_out[1] uo_out[1].n5 0.0730806
R1380 uo_out[3].n0 uo_out[3].t0 313.104
R1381 uo_out[3].t1 uo_out[3].n0 265.769
R1382 uo_out[3] uo_out[3].t1 262.318
R1383 uo_out[3].n2 uo_out[3] 19.5328
R1384 uo_out[3].n2 uo_out[3].n1 13.8005
R1385 uo_out[3].n1 uo_out[3].n0 7.17626
R1386 uo_out[3].n1 uo_out[3] 4.84898
R1387 uo_out[3] uo_out[3].n2 0.0529194
R1388 uo_out[2].n2 uo_out[2].t0 313.104
R1389 uo_out[2].n0 uo_out[2].t2 294.557
R1390 uo_out[2].t1 uo_out[2].n2 265.769
R1391 uo_out[2] uo_out[2].t1 262.318
R1392 uo_out[2].n0 uo_out[2].t3 211.01
R1393 uo_out[2].n1 uo_out[2].n0 152
R1394 uo_out[2].n5 uo_out[2] 16.2155
R1395 uo_out[2].n4 uo_out[2].n1 11.6311
R1396 uo_out[2].n4 uo_out[2].n3 9.3005
R1397 uo_out[2].n3 uo_out[2] 7.17626
R1398 uo_out[2].n3 uo_out[2].n2 4.84898
R1399 uo_out[2].n5 uo_out[2].n4 4.51042
R1400 uo_out[2].n1 uo_out[2] 1.37896
R1401 uo_out[2] uo_out[2].n5 0.0730806
C0 m2_15474_32386# m1_15474_32386# 2.03601f
C1 m4_10182_17306# m3_10182_17306# 47.1973f
C2 m1_18496_33616# m2_18496_33616# 2.03601f
C3 m1_4416_25486# m2_4416_25486# 2.03601f
C4 m1_20662_15338# m2_20662_15338# 2.03601f
C5 m2_7076_29088# m1_7076_29088# 2.03601f
C6 m2_22770_17310# m1_22770_17310# 2.03601f
C7 m1_22770_15390# m2_22770_15390# 2.03601f
C8 m1_3616_20266# m2_3616_20266# 2.03601f
C9 m1_21182_30146# m2_21182_30146# 2.03601f
C10 m3_11508_25704# m2_11508_25704# 71.142296f
C11 m1_24714_24800# m2_24714_24800# 2.03601f
C12 m1_7564_42050# m2_7564_42050# 2.03601f
C13 m1_14954_13098# m2_14954_13098# 2.03601f
C14 m1_4416_23566# m2_4416_23566# 2.03601f
C15 m1_15474_34306# m2_15474_34306# 2.03601f
C16 m2_14954_11178# m1_14954_11178# 2.03601f
C17 m2_10182_17306# m3_10182_17306# 48.4105f
C18 m2_12384_34074# m1_12384_34074# 2.03601f
C19 m2_10182_17306# m1_10182_17306# 75.185295f
C20 m2_5328_26928# m1_5328_26928# 2.03601f
C21 m1_6556_16396# m2_6556_16396# 2.03601f
C22 m1_24658_19894# m2_24658_19894# 2.03601f
C23 m1_6556_14476# m2_6556_14476# 2.03601f
C24 m3_11508_25704# m4_11508_25704# 69.3594f
C25 m1_24714_26720# m2_24714_26720# 2.03601f
C26 m1_18496_31696# m2_18496_31696# 2.03601f
C27 m1_25498_23336# m2_25498_23336# 2.03601f
C28 m2_12528_42110# m1_12528_42110# 2.03601f
C29 m1_11508_25704# m2_11508_25704# 0.11049p
C30 m1_7076_31008# m2_7076_31008# 2.03601f
C31 m2_11864_11410# m1_11864_11410# 2.03601f
C32 m1_5328_28848# m2_5328_28848# 2.03601f
C33 m1_4708_16904# m2_4708_16904# 2.03601f
C34 m1_8978_14462# m2_8978_14462# 2.03601f
C35 m1_3616_22186# m2_3616_22186# 2.03601f
C36 m2_9500_32942# m1_9500_32942# 2.03601f
C37 m1_24658_17974# m2_24658_17974# 2.03601f
C38 m2_4708_18824# m1_4708_18824# 2.03601f
C39 VDPWR VAPWR 21.118801f
C40 m1_11864_13330# m2_11864_13330# 2.03601f
C41 m1_9500_31022# m2_9500_31022# 2.03601f
C42 m1_8978_12542# m2_8978_12542# 2.03601f
C43 m2_23290_27874# m1_23290_27874# 2.03601f
C44 m1_10788_42050# m2_10788_42050# 2.03601f
C45 m1_17976_13788# m2_17976_13788# 2.03601f
C46 m1_21182_32066# m2_21182_32066# 2.03601f
C47 m2_17976_11868# m1_17976_11868# 2.03601f
C48 m1_23290_29794# m2_23290_29794# 2.03601f
C49 m1_25498_21416# m2_25498_21416# 2.03601f
C50 m1_12384_32154# m2_12384_32154# 2.03601f
C51 m2_9304_42110# m1_9304_42110# 2.03601f
C52 m2_20662_13418# m1_20662_13418# 2.03601f
C53 ua[0] VGND 29.2896f
C54 uo_out[0] VGND 3.93899f
C55 uo_out[3] VGND 1.88505f
C56 VAPWR VGND 0.142229p
C57 VDPWR VGND 51.147964f
C58 m4_10182_17306# VGND 9.38538f $ **FLOATING
C59 m4_11508_25704# VGND 7.22411f $ **FLOATING
C60 m3_10182_17306# VGND 10.656599f $ **FLOATING
C61 m3_11508_25704# VGND 8.43615f $ **FLOATING
C62 m2_10182_17306# VGND 9.82879f $ **FLOATING
C63 m2_11508_25704# VGND 7.81967f $ **FLOATING
C64 m1_10182_17306# VGND 25.3587f $ **FLOATING
C65 m1_11508_25704# VGND 30.364098f $ **FLOATING
C66 ring_0/skullfet_inverter_16.A VGND 4.7412f
C67 ring_0/skullfet_inverter_17.A VGND 4.82913f
C68 ring_0/skullfet_inverter_15.A VGND 4.9312f
C69 ring_0/skullfet_inverter_18.A VGND 4.98339f
C70 ring_0/skullfet_inverter_14.A VGND 5.03686f
C71 ring_0/skullfet_inverter_19.A VGND 4.79856f
C72 ring_0/skullfet_inverter_13.A VGND 4.80717f
C73 ring_0/skullfet_inverter_20.A VGND 4.93069f
C74 ring_0/skullfet_inverter_12.A VGND 6.09378f
C75 ring_0/skullfet_inverter_20.Y VGND 5.87716f
C76 ring_0/skullfet_inverter_11.A VGND 5.42552f
C77 ring_0/skullfet_inverter_1.A VGND 5.68048f
C78 ring_0/skullfet_inverter_10.A VGND 5.3549f
C79 ring_0/skullfet_inverter_2.A VGND 5.93378f
C80 ring_0/skullfet_inverter_9.A VGND 4.59492f
C81 ring_0/skullfet_inverter_3.A VGND 5.00062f
C82 ring_0/skullfet_inverter_4.A VGND 5.01468f
C83 ring_0/skullfet_inverter_7.A VGND 4.92037f
C84 ring_0/skullfet_inverter_6.A VGND 4.74003f
C85 ring_0/skullfet_inverter_5.A VGND 4.83065f
C86 skullfet_3v3_buffer.A VGND 12.652499f
C87 VDPWR.n3 VGND 7.05427f
C88 VAPWR.n67 VGND 2.60392f
C89 VAPWR.n69 VGND 16.1581f
.ends

