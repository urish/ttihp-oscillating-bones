magic
tech sky130A
magscale 1 2
timestamp 1735638153
<< metal1 >>
rect -586 10570 330 10670
rect 1764 10570 2596 10670
rect -3538 10338 -2760 10438
rect -1326 10434 -1126 10438
rect -586 10434 -486 10570
rect -1326 10338 -486 10434
rect -3538 9310 -3438 10338
rect -1220 10334 -486 10338
rect 2496 9980 2596 10570
rect 2496 9880 3352 9980
rect 4786 9880 5414 9980
rect -4090 9306 -3438 9310
rect -6170 9206 -5644 9306
rect -4210 9210 -3438 9306
rect -4210 9206 -4010 9210
rect -6170 7374 -6070 9206
rect 5314 8428 5414 9880
rect 5838 8428 6038 8430
rect 5314 8330 6038 8428
rect 7472 8330 7816 8430
rect 5314 8328 5906 8330
rect -6546 7372 -6070 7374
rect -8268 7272 -8068 7372
rect -6634 7274 -6070 7372
rect -6634 7272 -6434 7274
rect -8268 5212 -8168 7272
rect 7716 6158 7816 8330
rect 7716 6058 8146 6158
rect 9580 6058 9948 6158
rect -10016 5112 -9816 5212
rect -8382 5120 -8168 5212
rect -8382 5112 -8182 5120
rect -10016 3450 -9916 5112
rect 9848 4812 9948 6058
rect 9848 4712 11180 4812
rect -10016 3350 -9106 3450
rect -10994 1850 -10894 1864
rect -9206 1850 -9106 3350
rect 11080 3084 11180 4712
rect 9348 2984 9548 3084
rect 10982 2984 11182 3084
rect -10994 1750 -10728 1850
rect -9294 1750 -9094 1850
rect -10994 66 -10894 1750
rect -10994 -34 -9894 66
rect -9994 -1450 -9894 -34
rect 9348 -300 9448 2984
rect 9348 -400 10354 -300
rect 11788 -400 12170 -300
rect -11728 -1550 -11528 -1450
rect -10094 -1550 -9894 -1450
rect -11728 -3430 -11628 -1550
rect 12070 -1980 12170 -400
rect 11016 -2080 12170 -1980
rect -11728 -3530 -10922 -3430
rect -11022 -4804 -10922 -3530
rect 11016 -3764 11116 -2080
rect 9196 -3864 9500 -3764
rect 10934 -3864 11134 -3764
rect -11022 -4904 -10450 -4804
rect -9116 -4924 -8732 -4824
rect -8832 -7272 -8732 -4924
rect 9196 -6358 9296 -3864
rect 7244 -6458 7604 -6358
rect 9038 -6458 9296 -6358
rect -8832 -7372 -8610 -7272
rect -7176 -7276 -6976 -7272
rect -7176 -7372 -6514 -7276
rect -8832 -7376 -8732 -7372
rect -7096 -7376 -6514 -7372
rect -6614 -9206 -6514 -7376
rect 7244 -8328 7344 -6458
rect 9196 -6462 9296 -6458
rect 6968 -8330 7344 -8328
rect 5296 -8332 5496 -8330
rect 4810 -8430 5496 -8332
rect 6930 -8428 7344 -8330
rect 6930 -8430 7130 -8428
rect 4810 -8432 5374 -8430
rect -6632 -9306 -6188 -9206
rect -4754 -9210 -4554 -9206
rect -4754 -9306 -3900 -9210
rect -4656 -9310 -3900 -9306
rect -4000 -10338 -3900 -9310
rect 4810 -9880 4910 -8432
rect 1998 -9980 2810 -9880
rect 4244 -9980 4910 -9880
rect -1790 -10338 -932 -10334
rect -4000 -10438 -3302 -10338
rect -1868 -10434 -932 -10338
rect -1868 -10438 -1668 -10434
rect -1032 -10570 -932 -10434
rect -1032 -10670 -212 -10570
rect 1222 -10578 1422 -10570
rect 1998 -10578 2098 -9980
rect 1222 -10670 2098 -10578
rect 1318 -10678 2098 -10670
<< metal2 >>
rect -199 12870 200 12872
rect -359 12867 359 12870
rect -518 12862 518 12867
rect -677 12855 677 12862
rect -836 12846 836 12855
rect -995 12835 995 12846
rect -1154 12823 1154 12835
rect -1313 12808 1313 12823
rect -1471 12791 1471 12808
rect -1630 12772 1630 12791
rect -1788 12751 1788 12772
rect -1946 12728 1946 12751
rect -2103 12703 2103 12728
rect -2260 12676 2260 12703
rect -2417 12647 2417 12676
rect -2574 12616 2574 12647
rect -2730 12583 2730 12616
rect -2886 12549 2886 12583
rect -3041 12512 3041 12549
rect -3196 12473 3196 12512
rect -3351 12470 3351 12473
rect -3351 12467 -118 12470
rect 118 12467 3351 12470
rect -3351 12462 -277 12467
rect 277 12462 3351 12467
rect -3351 12455 -436 12462
rect 330 12455 3351 12462
rect -3351 12446 -595 12455
rect -3351 12435 -754 12446
rect -3351 12433 -913 12435
rect -3505 12423 -913 12433
rect -3505 12408 -1071 12423
rect -3505 12391 -1230 12408
rect 330 12407 467 12455
rect 595 12446 3351 12455
rect 754 12435 3351 12446
rect 913 12433 3351 12435
rect 913 12423 3505 12433
rect 1071 12408 3505 12423
rect -3505 12390 -1388 12391
rect -3658 12372 -1388 12390
rect -3658 12351 -1546 12372
rect -3658 12346 -1703 12351
rect -3811 12328 -1703 12346
rect -3811 12303 -1860 12328
rect -3811 12300 -2017 12303
rect -3964 12276 -2017 12300
rect -3964 12251 -2174 12276
rect -4115 12247 -2174 12251
rect -4115 12216 -2330 12247
rect -4115 12201 -2486 12216
rect -4266 12183 -2486 12201
rect -4266 12149 -2641 12183
rect -4417 12112 -2796 12149
rect -4417 12095 -2951 12112
rect -4567 12073 -2951 12095
rect -4567 12039 -3105 12073
rect -4716 12033 -3105 12039
rect -4716 11990 -3258 12033
rect -4716 11982 -3411 11990
rect -4864 11946 -3411 11982
rect -4864 11922 -3564 11946
rect -5012 11900 -3564 11922
rect -5012 11861 -3715 11900
rect -5159 11851 -3715 11861
rect -5159 11801 -3866 11851
rect -5159 11797 -4017 11801
rect -5305 11749 -4017 11797
rect -5305 11732 -4167 11749
rect -2760 11738 -2670 12149
rect 330 11970 420 12407
rect 1230 12391 3505 12408
rect 1388 12390 3505 12391
rect 1388 12372 3658 12390
rect 1546 12351 3658 12372
rect 1703 12346 3658 12351
rect 1703 12328 3811 12346
rect 1860 12303 3811 12328
rect 2017 12300 3811 12303
rect 2017 12276 3964 12300
rect 2174 12251 3964 12276
rect 2174 12247 4115 12251
rect 2330 12216 4115 12247
rect 2486 12201 4115 12216
rect 2486 12183 4266 12201
rect 2641 12149 4266 12183
rect 2796 12112 4417 12149
rect 2951 12095 4417 12112
rect 2951 12073 4567 12095
rect 3105 12039 4567 12073
rect 3105 12033 4716 12039
rect 3258 11990 4716 12033
rect 3352 11982 4716 11990
rect 3352 11946 4864 11982
rect -5450 11695 -4167 11732
rect -5450 11665 -4316 11695
rect -5595 11639 -4316 11665
rect -5595 11597 -4464 11639
rect -5739 11582 -4464 11597
rect -5739 11526 -4612 11582
rect -5881 11522 -4612 11526
rect -5881 11461 -4759 11522
rect -5881 11454 -4905 11461
rect -6023 11397 -4905 11454
rect -6023 11380 -5050 11397
rect -6164 11332 -5050 11380
rect -6164 11304 -5195 11332
rect -6304 11265 -5195 11304
rect 3352 11280 3442 11946
rect 3564 11922 4864 11946
rect 3564 11900 5012 11922
rect 3715 11861 5012 11900
rect 3715 11851 5159 11861
rect 3866 11801 5159 11851
rect 4017 11797 5159 11801
rect 4017 11749 5305 11797
rect 4167 11732 5305 11749
rect 4167 11695 5450 11732
rect 4316 11665 5450 11695
rect 4316 11639 5595 11665
rect 4464 11597 5595 11639
rect 4464 11582 5739 11597
rect 4612 11526 5739 11582
rect 4612 11522 5881 11526
rect 4759 11461 5881 11522
rect 4905 11454 5881 11461
rect 4905 11397 6023 11454
rect 5050 11380 6023 11397
rect 5050 11332 6164 11380
rect 5195 11304 6164 11332
rect 5195 11265 6304 11304
rect -6304 11226 -5339 11265
rect -6443 11197 -5339 11226
rect 5339 11226 6304 11265
rect 5339 11197 6443 11226
rect -6443 11147 -5481 11197
rect -6581 11126 -5481 11147
rect 5481 11147 6443 11197
rect 5481 11126 6581 11147
rect -6581 11066 -5554 11126
rect -6718 11054 -5554 11066
rect 5623 11066 6581 11126
rect 5623 11054 6718 11066
rect -6718 10983 -5764 11054
rect -6855 10980 -5764 10983
rect -6855 10904 -5904 10980
rect -6855 10899 -6043 10904
rect -6989 10826 -6043 10899
rect -6989 10813 -6181 10826
rect -7123 10747 -6181 10813
rect -7123 10725 -6318 10747
rect -7256 10666 -6318 10725
rect -7256 10635 -6455 10666
rect -7388 10583 -6455 10635
rect -5644 10606 -5554 11054
rect 5764 10983 6718 11054
rect 5764 10980 6855 10983
rect 5904 10904 6855 10980
rect 6038 10899 6855 10904
rect 6038 10826 6989 10899
rect -7388 10544 -6589 10583
rect -7519 10499 -6589 10544
rect -7519 10451 -6723 10499
rect -7648 10413 -6723 10451
rect -7648 10357 -6856 10413
rect -7776 10325 -6856 10357
rect -7776 10261 -6988 10325
rect -7903 10235 -6988 10261
rect -7903 10163 -7119 10235
rect -8029 10144 -7119 10163
rect -8029 10064 -7248 10144
rect -8154 10051 -7248 10064
rect -8154 9963 -7376 10051
rect -8277 9957 -7376 9963
rect -8277 9861 -7503 9957
rect -8399 9763 -7629 9861
rect -8399 9757 -7754 9763
rect -8520 9664 -7754 9757
rect 6038 9730 6128 10826
rect 6181 10813 6989 10826
rect 6181 10747 7123 10813
rect 6318 10725 7123 10747
rect 6318 10666 7256 10725
rect 6455 10635 7256 10666
rect 6455 10583 7388 10635
rect 6589 10544 7388 10583
rect 6589 10499 7519 10544
rect 6723 10451 7519 10499
rect 6723 10413 7648 10451
rect 6856 10357 7648 10413
rect 6856 10325 7776 10357
rect 6988 10261 7776 10325
rect 6988 10235 7903 10261
rect 7119 10163 7903 10235
rect 7119 10144 8029 10163
rect 7248 10064 8029 10144
rect 7248 10051 8154 10064
rect 7376 9963 8154 10051
rect 7376 9957 8277 9963
rect 7503 9861 8277 9957
rect 7629 9763 8399 9861
rect 7754 9757 8399 9763
rect 7754 9664 8520 9757
rect -8520 9652 -7877 9664
rect -8639 9563 -7877 9652
rect 7877 9652 8520 9664
rect 7877 9563 8639 9652
rect -8639 9545 -7999 9563
rect -8757 9461 -7999 9545
rect 7999 9545 8639 9563
rect 7999 9461 8757 9545
rect -8757 9437 -8120 9461
rect -8874 9357 -8120 9437
rect 8120 9437 8757 9461
rect 8120 9357 8874 9437
rect -8874 9327 -8239 9357
rect -8989 9252 -8239 9327
rect 8239 9327 8874 9357
rect 8239 9252 8989 9327
rect -8989 9216 -8357 9252
rect -9103 9145 -8357 9216
rect 8357 9216 8989 9252
rect -9103 9103 -8474 9145
rect -9216 9037 -8474 9103
rect -9216 8989 -8589 9037
rect -9327 8927 -8589 8989
rect -9327 8874 -8703 8927
rect -9437 8872 -8703 8874
rect -9437 8782 -7978 8872
rect -9437 8757 -8816 8782
rect -9545 8703 -8816 8757
rect -9545 8639 -8927 8703
rect -8068 8672 -7978 8782
rect -9652 8589 -8927 8639
rect -9652 8520 -9037 8589
rect -9757 8474 -9037 8520
rect -9757 8399 -9145 8474
rect -9861 8357 -9145 8399
rect -9861 8277 -9252 8357
rect -9963 8239 -9252 8277
rect -2760 8259 -2670 8938
rect -199 8598 200 8600
rect 330 8598 420 9170
rect 8357 9145 9103 9216
rect 8474 9103 9103 9145
rect 8474 9037 9216 9103
rect 8589 8989 9216 9037
rect 8589 8927 9327 8989
rect 8703 8874 9327 8927
rect 8703 8816 9437 8874
rect 8816 8757 9437 8816
rect 8816 8703 9545 8757
rect -346 8594 420 8598
rect 8927 8639 9545 8703
rect -493 8588 493 8594
rect 8927 8589 9652 8639
rect -639 8579 639 8588
rect -785 8568 785 8579
rect -932 8553 932 8568
rect -1078 8537 1078 8553
rect -1223 8518 1223 8537
rect 9037 8520 9652 8589
rect -1369 8496 1369 8518
rect -1514 8472 1514 8496
rect -1658 8445 1658 8472
rect -1802 8416 1802 8445
rect -1946 8384 1946 8416
rect -2089 8350 2089 8384
rect -2232 8313 2232 8350
rect -2374 8274 2374 8313
rect -9963 8154 -9357 8239
rect -2760 8232 -2619 8259
rect -2515 8232 2515 8274
rect -2760 8198 2655 8232
rect -2760 8194 -93 8198
rect 93 8194 2655 8198
rect -2760 8188 -239 8194
rect 239 8188 2655 8194
rect -10064 8120 -9357 8154
rect -2795 8179 -385 8188
rect 385 8179 2795 8188
rect -2795 8168 -532 8179
rect 532 8168 2795 8179
rect -2795 8153 -678 8168
rect 678 8153 2795 8168
rect -2795 8142 -823 8153
rect -2934 8137 -823 8142
rect 823 8142 2795 8153
rect 823 8137 2934 8142
rect -10064 8029 -9461 8120
rect -2934 8118 -969 8137
rect 969 8118 2934 8137
rect -2934 8096 -1114 8118
rect 1114 8096 2934 8118
rect -2934 8093 -1258 8096
rect -3072 8072 -1258 8093
rect 1258 8093 2934 8096
rect 1258 8072 3072 8093
rect -3072 8045 -1402 8072
rect 1402 8045 3072 8072
rect -3072 8042 -1546 8045
rect -10163 7999 -9461 8029
rect -3210 8016 -1546 8042
rect 1546 8042 3072 8045
rect 1546 8016 3210 8042
rect -10163 7903 -9563 7999
rect -3210 7988 -1689 8016
rect -3346 7984 -1689 7988
rect 1689 7988 3210 8016
rect 3352 8005 3442 8480
rect 9037 8474 9757 8520
rect 9145 8399 9757 8474
rect 9145 8357 9861 8399
rect 9252 8277 9861 8357
rect 9252 8239 9963 8277
rect 9357 8154 9963 8239
rect 9357 8120 10064 8154
rect 9461 8029 10064 8120
rect 9461 8005 10163 8029
rect 3285 7988 3442 8005
rect 1689 7984 3442 7988
rect -3346 7950 -1832 7984
rect 1832 7950 3442 7984
rect -3346 7932 -1974 7950
rect -10261 7877 -9563 7903
rect -3482 7913 -1974 7932
rect 1974 7932 3442 7950
rect 1974 7913 3482 7932
rect -10261 7776 -9664 7877
rect -3482 7874 -2115 7913
rect 2115 7874 3482 7913
rect -3482 7873 -2255 7874
rect -3616 7832 -2255 7873
rect 2255 7873 3482 7874
rect 8146 7915 10163 8005
rect 2255 7832 3616 7873
rect -3616 7812 -2395 7832
rect -10357 7754 -9664 7776
rect -10357 7648 -9763 7754
rect -10451 7629 -9763 7648
rect -10451 7519 -9861 7629
rect -10544 7503 -9861 7519
rect -10544 7388 -9957 7503
rect -10635 7376 -9957 7388
rect -10635 7256 -10051 7376
rect -10725 7248 -10051 7256
rect -10725 7123 -10144 7248
rect -10813 7119 -10144 7123
rect -10813 6989 -10235 7119
rect -10899 6988 -10235 6989
rect -10899 6856 -10325 6988
rect -10899 6855 -10413 6856
rect -10983 6723 -10413 6855
rect -10983 6718 -10499 6723
rect -11066 6645 -10499 6718
rect -11066 6581 -9726 6645
rect -11147 6555 -9726 6581
rect -11147 6455 -10583 6555
rect -9816 6512 -9726 6555
rect -5644 6634 -5554 7806
rect -3749 7788 -2395 7812
rect 2395 7812 3616 7832
rect 2395 7788 3749 7812
rect -3749 7749 -2534 7788
rect -3882 7742 -2534 7749
rect 2534 7749 3749 7788
rect 2534 7742 3882 7749
rect -3882 7693 -2672 7742
rect 2672 7693 3882 7742
rect -3882 7684 -2810 7693
rect -4013 7642 -2810 7684
rect 2810 7684 3882 7693
rect 2810 7642 4013 7684
rect -4013 7616 -2946 7642
rect -4143 7588 -2946 7616
rect 2946 7616 4013 7642
rect 2946 7588 4143 7616
rect -4143 7546 -3082 7588
rect -4272 7532 -3082 7546
rect 3082 7546 4143 7588
rect 3082 7532 4272 7546
rect -4272 7474 -3216 7532
rect -4399 7473 -3216 7474
rect 3216 7474 4272 7532
rect 3216 7473 4400 7474
rect -4399 7412 -3349 7473
rect 3349 7412 4400 7473
rect 8146 7458 8236 7915
rect 9563 7903 10163 7915
rect 9563 7877 10261 7903
rect 9664 7776 10261 7877
rect 9664 7754 10357 7776
rect 9763 7648 10357 7754
rect 9763 7629 10451 7648
rect 9861 7519 10451 7629
rect 9861 7503 10544 7519
rect -4399 7400 -3482 7412
rect -4526 7349 -3482 7400
rect 3482 7400 4400 7412
rect 3482 7349 4526 7400
rect 9957 7388 10544 7503
rect 9957 7376 10635 7388
rect -4526 7323 -3613 7349
rect -4651 7284 -3613 7323
rect 3613 7323 4526 7349
rect 3613 7284 4651 7323
rect -4651 7244 -3743 7284
rect -4774 7216 -3743 7244
rect 3743 7244 4651 7284
rect 10051 7256 10635 7376
rect 10051 7248 10725 7256
rect 3743 7216 4774 7244
rect -4774 7163 -3872 7216
rect -4897 7146 -3872 7163
rect 3872 7163 4774 7216
rect 3872 7146 4897 7163
rect -4897 7080 -3999 7146
rect -5018 7074 -3999 7080
rect 4000 7080 4897 7146
rect 10144 7123 10725 7248
rect 10144 7119 10813 7123
rect 4000 7074 5018 7080
rect -5018 7000 -4126 7074
rect 4126 7000 5018 7074
rect -5018 6995 -4251 7000
rect -5137 6923 -4251 6995
rect 4251 6995 5018 7000
rect 4251 6923 5137 6995
rect 10235 6989 10813 7119
rect 10235 6988 10899 6989
rect -5137 6908 -4374 6923
rect -5255 6844 -4374 6908
rect 4374 6908 5137 6923
rect 4374 6844 5255 6908
rect -5255 6819 -4497 6844
rect -5371 6763 -4497 6819
rect 4497 6819 5255 6844
rect 4497 6773 5371 6819
rect 6038 6773 6128 6930
rect 10325 6856 10899 6988
rect 4497 6763 6128 6773
rect -5371 6728 -4618 6763
rect -5486 6680 -4618 6728
rect 4618 6683 6128 6763
rect 10413 6855 10899 6856
rect 10413 6723 10983 6855
rect 10499 6718 10983 6723
rect 4618 6680 5486 6683
rect -5486 6634 -4737 6680
rect -5644 6595 -4737 6634
rect 4737 6634 5486 6680
rect 4737 6595 5599 6634
rect -5644 6539 -4855 6595
rect -5710 6508 -4855 6539
rect 4855 6539 5599 6595
rect 10499 6589 11066 6718
rect 10583 6581 11066 6589
rect 4855 6508 5710 6539
rect -11147 6443 -10666 6455
rect -11226 6318 -10666 6443
rect -5710 6442 -4971 6508
rect -5820 6419 -4971 6442
rect 4971 6442 5710 6508
rect 10583 6455 11147 6581
rect 10666 6443 11147 6455
rect 4971 6419 5820 6442
rect -5820 6343 -5086 6419
rect -5928 6328 -5086 6343
rect 5086 6343 5820 6419
rect 5086 6328 5928 6343
rect -11226 6304 -10747 6318
rect -11304 6181 -10747 6304
rect -5928 6242 -5199 6328
rect -6035 6234 -5199 6242
rect 5199 6242 5928 6328
rect 10666 6318 11226 6443
rect 10747 6304 11226 6318
rect 5199 6234 6035 6242
rect -11304 6164 -10826 6181
rect -11380 6043 -10826 6164
rect -6035 6139 -5310 6234
rect 5310 6139 6035 6234
rect 10747 6181 11304 6304
rect 10826 6164 11304 6181
rect -11380 6023 -10904 6043
rect -6139 6042 -5420 6139
rect 5420 6042 6139 6139
rect 10826 6043 11380 6164
rect -6139 6035 -5528 6042
rect -11454 5904 -10904 6023
rect -6242 5943 -5528 6035
rect 5528 6035 6139 6042
rect 5528 5943 6242 6035
rect -6242 5928 -5635 5943
rect -11454 5881 -10980 5904
rect -11526 5764 -10980 5881
rect -8068 5765 -7978 5872
rect -6343 5842 -5635 5928
rect 5635 5928 6242 5943
rect 10904 6023 11380 6043
rect 5635 5842 6343 5928
rect 10904 5904 11454 6023
rect -6343 5820 -5739 5842
rect -6442 5765 -5739 5820
rect -11526 5739 -11054 5764
rect -11597 5623 -11054 5739
rect -8068 5739 -5739 5765
rect 5739 5820 6343 5842
rect 10980 5881 11454 5904
rect 5739 5739 6442 5820
rect 10980 5764 11526 5881
rect -8068 5675 -5842 5739
rect -8068 5672 -7978 5675
rect -6539 5635 -5842 5675
rect 5842 5710 6442 5739
rect 11054 5739 11526 5764
rect 5842 5635 6539 5710
rect -11597 5595 -11126 5623
rect -6539 5599 -5943 5635
rect -11665 5481 -11126 5595
rect -6634 5528 -5943 5599
rect 5943 5599 6539 5635
rect 11054 5623 11597 5739
rect 5943 5528 6634 5599
rect -6634 5486 -6042 5528
rect -11665 5450 -11197 5481
rect -11732 5339 -11197 5450
rect -6728 5420 -6042 5486
rect 6042 5486 6634 5528
rect 11126 5595 11597 5623
rect 6042 5420 6728 5486
rect 11126 5481 11665 5595
rect -6728 5371 -6139 5420
rect -11732 5305 -11265 5339
rect -11797 5195 -11265 5305
rect -6819 5310 -6139 5371
rect 6139 5371 6728 5420
rect 11197 5450 11665 5481
rect 6139 5310 6819 5371
rect 11197 5339 11732 5450
rect -6819 5255 -6234 5310
rect -6908 5199 -6234 5255
rect 6234 5255 6819 5310
rect 11265 5305 11732 5339
rect 6234 5199 6908 5255
rect -11797 5159 -11332 5195
rect -11861 5050 -11332 5159
rect -6908 5137 -6328 5199
rect -6995 5086 -6328 5137
rect 6328 5137 6908 5199
rect 11265 5195 11797 5305
rect 11332 5159 11797 5195
rect 6328 5086 6995 5137
rect -11861 5012 -11397 5050
rect -6995 5018 -6419 5086
rect -11922 4905 -11397 5012
rect -7080 4971 -6419 5018
rect 6419 5018 6995 5086
rect 11332 5050 11861 5159
rect 6419 4971 7080 5018
rect -11922 4864 -11461 4905
rect -7080 4897 -6508 4971
rect -11982 4759 -11461 4864
rect -7163 4855 -6508 4897
rect 6508 4897 7080 4971
rect 11397 5012 11861 5050
rect 11397 4905 11922 5012
rect 6508 4855 7163 4897
rect -7163 4774 -6595 4855
rect -11982 4716 -11522 4759
rect -12039 4612 -11522 4716
rect -7244 4737 -6595 4774
rect 6595 4774 7163 4855
rect 11461 4864 11922 4905
rect 6595 4737 7244 4774
rect 11461 4759 11982 4864
rect -7244 4651 -6680 4737
rect -7323 4618 -6680 4651
rect 6680 4651 7244 4737
rect 11522 4716 11982 4759
rect 6680 4618 7323 4651
rect -12039 4567 -11582 4612
rect -12095 4464 -11582 4567
rect -7323 4526 -6763 4618
rect -7400 4497 -6763 4526
rect 6763 4548 7323 4618
rect 8146 4548 8236 4658
rect 11522 4612 12039 4716
rect 11582 4584 12039 4612
rect 6763 4497 8236 4548
rect -12095 4417 -11639 4464
rect -12149 4316 -11639 4417
rect -7400 4399 -6844 4497
rect -7474 4374 -6844 4399
rect 6844 4458 8236 4497
rect 10892 4567 12039 4584
rect 10892 4494 12095 4567
rect 6844 4399 7400 4458
rect 6844 4374 7474 4399
rect 10892 4384 10982 4494
rect 11582 4464 12095 4494
rect 11639 4417 12095 4464
rect -12149 4266 -11695 4316
rect -7474 4272 -6923 4374
rect -12201 4167 -11695 4266
rect -7546 4251 -6923 4272
rect 6923 4272 7474 4374
rect 11639 4316 12149 4417
rect 6923 4251 7546 4272
rect -12201 4115 -11749 4167
rect -7546 4143 -7000 4251
rect -12251 4017 -11749 4115
rect -7616 4126 -7000 4143
rect 7000 4143 7546 4251
rect 11695 4266 12149 4316
rect 11695 4167 12201 4266
rect 7000 4126 7616 4143
rect -12251 3964 -11801 4017
rect -7616 4013 -7074 4126
rect -12300 3866 -11801 3964
rect -7684 3999 -7074 4013
rect 7074 4013 7616 4126
rect 11749 4115 12201 4167
rect 11749 4017 12251 4115
rect 7074 3999 7684 4013
rect -7684 3882 -7146 3999
rect -7749 3872 -7146 3882
rect 7146 3882 7684 3999
rect 11801 3964 12251 4017
rect 7146 3872 7749 3882
rect -12300 3811 -11851 3866
rect -12346 3715 -11851 3811
rect -7749 3749 -7216 3872
rect -7812 3743 -7216 3749
rect 7216 3749 7749 3872
rect 11801 3866 12300 3964
rect 11851 3811 12300 3866
rect 7216 3743 7812 3749
rect -12346 3658 -11900 3715
rect -12390 3564 -11900 3658
rect -9816 3602 -9726 3712
rect -7812 3616 -7284 3743
rect -7873 3613 -7284 3616
rect 7284 3616 7812 3743
rect 11851 3715 12346 3811
rect 11900 3658 12346 3715
rect 7284 3613 7873 3616
rect -7873 3602 -7349 3613
rect -12390 3505 -11946 3564
rect -9816 3512 -7349 3602
rect -12433 3411 -11946 3505
rect -7873 3482 -7349 3512
rect 7349 3482 7873 3613
rect 11900 3564 12390 3658
rect 11946 3505 12390 3564
rect -12433 3351 -11990 3411
rect -12473 3350 -11990 3351
rect -12473 3260 -10638 3350
rect -7932 3349 -7412 3482
rect 7412 3349 7932 3482
rect 11946 3411 12433 3505
rect -7932 3346 -7473 3349
rect -12473 3258 -11990 3260
rect -12473 3196 -12033 3258
rect -12512 3105 -12033 3196
rect -10728 3150 -10638 3260
rect -7988 3216 -7473 3346
rect 7473 3346 7932 3349
rect 11990 3351 12433 3411
rect 7473 3216 7988 3346
rect 11990 3258 12473 3351
rect -7988 3210 -7532 3216
rect -12512 3041 -12073 3105
rect -8042 3082 -7532 3210
rect 7532 3210 7988 3216
rect 7532 3082 8042 3210
rect 12033 3196 12473 3258
rect 12033 3105 12512 3196
rect -8042 3072 -7588 3082
rect -12549 2951 -12073 3041
rect -12549 2886 -12112 2951
rect -8093 2946 -7588 3072
rect 7588 3072 8042 3082
rect 7588 2946 8093 3072
rect 12073 3041 12512 3105
rect 12073 2951 12549 3041
rect -8093 2934 -7642 2946
rect -12583 2796 -12112 2886
rect -8142 2810 -7642 2934
rect 7642 2934 8093 2946
rect 7642 2810 8142 2934
rect -12583 2730 -12149 2796
rect -8142 2795 -7693 2810
rect -12616 2641 -12149 2730
rect -8188 2672 -7693 2795
rect 7693 2795 8142 2810
rect 12112 2886 12549 2951
rect 12112 2796 12583 2886
rect 7693 2672 8188 2795
rect -8188 2655 -7742 2672
rect -12616 2574 -12183 2641
rect -12647 2486 -12183 2574
rect -8232 2534 -7742 2655
rect 7742 2655 8188 2672
rect 12149 2730 12583 2796
rect 7742 2534 8232 2655
rect 12149 2641 12616 2730
rect -8232 2515 -7788 2534
rect -12647 2417 -12216 2486
rect -12676 2330 -12216 2417
rect -8274 2395 -7788 2515
rect 7788 2515 8232 2534
rect 12183 2574 12616 2641
rect 7788 2395 8274 2515
rect 12183 2486 12647 2574
rect -8274 2374 -7832 2395
rect -12676 2260 -12247 2330
rect -12703 2174 -12247 2260
rect -8313 2255 -7832 2374
rect 7832 2374 8274 2395
rect 12216 2417 12647 2486
rect 7832 2255 8313 2374
rect 12216 2330 12676 2417
rect -8313 2232 -7874 2255
rect -12703 2103 -12276 2174
rect -12728 2017 -12276 2103
rect -8350 2115 -7874 2232
rect 7874 2232 8313 2255
rect 12247 2260 12676 2330
rect 7874 2115 8350 2232
rect 12247 2174 12703 2260
rect -8350 2089 -7913 2115
rect -12728 1946 -12303 2017
rect -8384 1974 -7913 2089
rect 7913 2089 8350 2115
rect 12276 2103 12703 2174
rect 7913 1974 8384 2089
rect 12276 2017 12728 2103
rect -8384 1946 -7950 1974
rect -12751 1860 -12303 1946
rect -12751 1788 -12328 1860
rect -8416 1832 -7950 1946
rect 7950 1946 8384 1974
rect 12303 1946 12728 2017
rect 7950 1832 8416 1946
rect 12303 1860 12751 1946
rect -8416 1802 -7984 1832
rect -12772 1703 -12328 1788
rect -12772 1630 -12351 1703
rect -8445 1689 -7984 1802
rect 7984 1802 8416 1832
rect 7984 1689 8445 1802
rect 12328 1788 12751 1860
rect 12328 1703 12772 1788
rect -8445 1658 -8016 1689
rect -12791 1546 -12351 1630
rect -8472 1546 -8016 1658
rect 8016 1658 8445 1689
rect 8016 1546 8472 1658
rect 12351 1630 12772 1703
rect -12791 1471 -12372 1546
rect -8472 1514 -8045 1546
rect -12808 1388 -12372 1471
rect -8496 1402 -8045 1514
rect 8045 1514 8472 1546
rect 8045 1474 8496 1514
rect 10892 1474 10982 1584
rect 12351 1546 12791 1630
rect 8045 1402 10982 1474
rect -12808 1313 -12391 1388
rect -8496 1369 -8072 1402
rect -12823 1230 -12391 1313
rect -8518 1258 -8072 1369
rect 8072 1384 10982 1402
rect 12372 1471 12791 1546
rect 12372 1388 12808 1471
rect 8072 1307 8547 1384
rect 12391 1313 12808 1388
rect 8072 1258 8518 1307
rect -12823 1154 -12408 1230
rect -8518 1223 -8096 1258
rect -12835 1071 -12408 1154
rect -8537 1114 -8096 1223
rect 8096 1223 8518 1258
rect 12391 1230 12823 1313
rect 8096 1114 8537 1223
rect -8537 1078 -8118 1114
rect -12835 995 -12423 1071
rect -12846 913 -12423 995
rect -8553 969 -8118 1078
rect 8118 1078 8537 1114
rect 10354 1154 12823 1230
rect 10354 1140 12835 1154
rect 8118 969 8553 1078
rect 10354 1000 10444 1140
rect 12408 1071 12835 1140
rect -8553 932 -8137 969
rect -12846 836 -12435 913
rect -12855 754 -12435 836
rect -8568 823 -8137 932
rect 8137 932 8553 969
rect 12423 995 12835 1071
rect 8137 823 8568 932
rect 12423 913 12846 995
rect -8568 785 -8153 823
rect -12855 677 -12446 754
rect -12862 595 -12446 677
rect -8579 678 -8153 785
rect 8153 785 8568 823
rect 12435 836 12846 913
rect 8153 678 8579 785
rect 12435 754 12855 836
rect -8579 639 -8168 678
rect -12862 518 -12455 595
rect -12867 436 -12455 518
rect -8588 532 -8168 639
rect 8168 639 8579 678
rect 12446 677 12855 754
rect 8168 532 8588 639
rect 12446 595 12862 677
rect -8588 493 -8179 532
rect -12867 359 -12462 436
rect -12870 277 -12462 359
rect -8594 385 -8179 493
rect 8179 493 8588 532
rect 12455 518 12862 595
rect 8179 385 8594 493
rect 12455 436 12867 518
rect -12870 200 -12467 277
rect -12872 118 -12467 200
rect -10728 240 -10638 350
rect -8594 346 -8188 385
rect -8598 240 -8188 346
rect -10728 239 -8188 240
rect 8188 346 8594 385
rect 12462 359 12867 436
rect 8188 239 8598 346
rect 12462 277 12870 359
rect -10728 150 -8194 239
rect -12872 50 -12470 118
rect -8600 93 -8194 150
rect 8194 200 8598 239
rect 12467 200 12870 277
rect 8194 93 8600 200
rect 12467 118 12872 200
rect -12872 -40 -11438 50
rect -12872 -118 -12470 -40
rect -12872 -199 -12467 -118
rect -11528 -150 -11438 -40
rect -8600 -93 -8198 93
rect 8198 -93 8600 93
rect -8600 -199 -8194 -93
rect -12870 -277 -12467 -199
rect -8598 -239 -8194 -199
rect 8194 -200 8600 -93
rect 12470 -118 12872 118
rect 12467 -200 12872 -118
rect 8194 -239 8598 -200
rect -12870 -359 -12462 -277
rect -8598 -346 -8188 -239
rect -12867 -436 -12462 -359
rect -8594 -385 -8188 -346
rect 8188 -346 8598 -239
rect 12467 -277 12870 -200
rect 8188 -385 8594 -346
rect -12867 -518 -12455 -436
rect -8594 -493 -8179 -385
rect -12862 -595 -12455 -518
rect -8588 -532 -8179 -493
rect 8179 -493 8594 -385
rect 12462 -359 12870 -277
rect 12462 -436 12867 -359
rect 8179 -532 8588 -493
rect -12862 -677 -12446 -595
rect -8588 -639 -8168 -532
rect -12855 -754 -12446 -677
rect -8579 -678 -8168 -639
rect 8168 -639 8588 -532
rect 12455 -518 12867 -436
rect 12455 -595 12862 -518
rect 8168 -678 8579 -639
rect -12855 -836 -12435 -754
rect -8579 -785 -8153 -678
rect -12846 -913 -12435 -836
rect -8568 -823 -8153 -785
rect 8153 -785 8579 -678
rect 12446 -677 12862 -595
rect 12446 -754 12855 -677
rect 8153 -823 8568 -785
rect -12846 -995 -12423 -913
rect -8568 -932 -8137 -823
rect -12835 -1071 -12423 -995
rect -8553 -969 -8137 -932
rect 8137 -932 8568 -823
rect 12435 -836 12855 -754
rect 12435 -913 12846 -836
rect 8137 -969 8553 -932
rect -12835 -1154 -12408 -1071
rect -8553 -1078 -8118 -969
rect -12823 -1230 -12408 -1154
rect -8537 -1114 -8118 -1078
rect 8118 -1078 8553 -969
rect 12423 -995 12846 -913
rect 12423 -1071 12835 -995
rect 8118 -1114 8537 -1078
rect -8537 -1223 -8096 -1114
rect -12823 -1313 -12391 -1230
rect -12808 -1388 -12391 -1313
rect -8518 -1258 -8096 -1223
rect 8096 -1223 8537 -1114
rect 12408 -1154 12835 -1071
rect 8096 -1258 8518 -1223
rect 12408 -1230 12823 -1154
rect -8518 -1369 -8072 -1258
rect -12808 -1471 -12372 -1388
rect -12791 -1546 -12372 -1471
rect -8496 -1402 -8072 -1369
rect 8072 -1369 8518 -1258
rect 12391 -1313 12823 -1230
rect 8072 -1402 8496 -1369
rect 12391 -1388 12808 -1313
rect -8496 -1514 -8045 -1402
rect -8472 -1546 -8045 -1514
rect 8045 -1514 8496 -1402
rect 12372 -1471 12808 -1388
rect 8045 -1546 8472 -1514
rect 12372 -1546 12791 -1471
rect -12791 -1630 -12351 -1546
rect -12772 -1703 -12351 -1630
rect -8472 -1658 -8016 -1546
rect -8445 -1689 -8016 -1658
rect 8016 -1658 8472 -1546
rect 12351 -1630 12791 -1546
rect 8016 -1689 8445 -1658
rect -12772 -1788 -12328 -1703
rect -12751 -1860 -12328 -1788
rect -8445 -1802 -7984 -1689
rect -8416 -1832 -7984 -1802
rect 7984 -1802 8445 -1689
rect 12351 -1703 12772 -1630
rect 12328 -1788 12772 -1703
rect 7984 -1832 8416 -1802
rect -12751 -1946 -12303 -1860
rect -8416 -1946 -7950 -1832
rect -12728 -2017 -12303 -1946
rect -8384 -1974 -7950 -1946
rect 7950 -1910 8416 -1832
rect 10354 -1909 10444 -1800
rect 12328 -1860 12751 -1788
rect 10223 -1910 10934 -1909
rect 7950 -1974 10934 -1910
rect -12728 -2103 -12276 -2017
rect -8384 -2089 -7913 -1974
rect -12703 -2174 -12276 -2103
rect -8350 -2115 -7913 -2089
rect 7913 -1999 10934 -1974
rect 7913 -2000 10444 -1999
rect 7913 -2089 8384 -2000
rect 7913 -2115 8350 -2089
rect -12703 -2260 -12247 -2174
rect -8350 -2232 -7874 -2115
rect -12676 -2330 -12247 -2260
rect -8313 -2255 -7874 -2232
rect 7874 -2232 8350 -2115
rect 7874 -2255 8313 -2232
rect -12676 -2417 -12216 -2330
rect -8313 -2374 -7832 -2255
rect -12647 -2486 -12216 -2417
rect -8274 -2395 -7832 -2374
rect 7832 -2374 8313 -2255
rect 7832 -2395 8274 -2374
rect -12647 -2574 -12183 -2486
rect -8274 -2515 -7788 -2395
rect -12616 -2641 -12183 -2574
rect -8232 -2534 -7788 -2515
rect 7788 -2515 8274 -2395
rect 10844 -2464 10934 -1999
rect 12303 -1946 12751 -1860
rect 12303 -2017 12728 -1946
rect 12276 -2103 12728 -2017
rect 12276 -2174 12703 -2103
rect 12247 -2260 12703 -2174
rect 12247 -2330 12676 -2260
rect 12216 -2417 12676 -2330
rect 12216 -2486 12647 -2417
rect 7788 -2534 8232 -2515
rect -12616 -2730 -12149 -2641
rect -8232 -2655 -7742 -2534
rect -12583 -2796 -12149 -2730
rect -8188 -2672 -7742 -2655
rect 7742 -2655 8232 -2534
rect 12183 -2574 12647 -2486
rect 12183 -2641 12616 -2574
rect 7742 -2672 8188 -2655
rect -8188 -2795 -7693 -2672
rect -12583 -2886 -12112 -2796
rect -12549 -2951 -12112 -2886
rect -8142 -2810 -7693 -2795
rect 7693 -2795 8188 -2672
rect 12149 -2730 12616 -2641
rect 7693 -2810 8142 -2795
rect 12149 -2796 12583 -2730
rect -8142 -2934 -7642 -2810
rect -8093 -2946 -7642 -2934
rect 7642 -2934 8142 -2810
rect 12112 -2886 12583 -2796
rect 7642 -2946 8093 -2934
rect -12549 -3041 -12073 -2951
rect -12512 -3105 -12073 -3041
rect -11528 -3059 -11438 -2950
rect -8093 -3059 -7588 -2946
rect -11528 -3082 -7588 -3059
rect 7588 -3072 8093 -2946
rect 12112 -2951 12549 -2886
rect 12073 -3041 12549 -2951
rect 7588 -3082 8042 -3072
rect -12512 -3196 -12033 -3105
rect -11528 -3149 -7532 -3082
rect -11528 -3150 -11438 -3149
rect -12473 -3258 -12033 -3196
rect -8042 -3210 -7532 -3149
rect -7988 -3216 -7532 -3210
rect 7532 -3210 8042 -3082
rect 12073 -3105 12512 -3041
rect 12033 -3196 12512 -3105
rect 7532 -3216 7988 -3210
rect -12473 -3287 -11990 -3258
rect -12473 -3351 -9024 -3287
rect -7988 -3346 -7473 -3216
rect -12433 -3377 -9024 -3351
rect -12433 -3411 -11990 -3377
rect -12433 -3505 -11946 -3411
rect -12390 -3564 -11946 -3505
rect -9114 -3514 -9024 -3377
rect -7932 -3349 -7473 -3346
rect 7473 -3346 7988 -3216
rect 12033 -3258 12473 -3196
rect 7473 -3349 7932 -3346
rect -7932 -3482 -7412 -3349
rect 7412 -3482 7932 -3349
rect 11990 -3351 12473 -3258
rect 11990 -3411 12433 -3351
rect -12390 -3658 -11900 -3564
rect -7873 -3613 -7349 -3482
rect 7349 -3613 7873 -3482
rect 11946 -3505 12433 -3411
rect 11946 -3564 12390 -3505
rect -7873 -3616 -7284 -3613
rect -12346 -3715 -11900 -3658
rect -12346 -3811 -11851 -3715
rect -7812 -3743 -7284 -3616
rect 7284 -3616 7873 -3613
rect 7284 -3743 7812 -3616
rect 11900 -3658 12390 -3564
rect 11900 -3715 12346 -3658
rect -7812 -3749 -7216 -3743
rect -12300 -3866 -11851 -3811
rect -12300 -3964 -11801 -3866
rect -7749 -3872 -7216 -3749
rect 7216 -3749 7812 -3743
rect 7216 -3872 7749 -3749
rect 11851 -3811 12346 -3715
rect 11851 -3866 12300 -3811
rect -7749 -3882 -7146 -3872
rect -12251 -4017 -11801 -3964
rect -7684 -4000 -7146 -3882
rect 7146 -3882 7749 -3872
rect 7146 -4000 7684 -3882
rect -7684 -4013 -7074 -4000
rect -12251 -4115 -11749 -4017
rect -12201 -4167 -11749 -4115
rect -7616 -4126 -7074 -4013
rect 7074 -4013 7684 -4000
rect 11801 -3964 12300 -3866
rect 7074 -4126 7616 -4013
rect 11801 -4017 12251 -3964
rect -7616 -4143 -7000 -4126
rect -12201 -4266 -11695 -4167
rect -12149 -4316 -11695 -4266
rect -7546 -4251 -7000 -4143
rect 7000 -4143 7616 -4126
rect 11749 -4115 12251 -4017
rect 7000 -4251 7546 -4143
rect 11749 -4167 12201 -4115
rect -7546 -4272 -6923 -4251
rect -12149 -4417 -11639 -4316
rect -7474 -4374 -6923 -4272
rect 6923 -4272 7546 -4251
rect 11695 -4266 12201 -4167
rect 6923 -4374 7474 -4272
rect 11695 -4316 12149 -4266
rect -7474 -4400 -6844 -4374
rect -12095 -4464 -11639 -4417
rect -12095 -4567 -11582 -4464
rect -7400 -4497 -6844 -4400
rect 6844 -4400 7474 -4374
rect 6844 -4497 7400 -4400
rect 11639 -4417 12149 -4316
rect 11639 -4464 12095 -4417
rect -7400 -4526 -6763 -4497
rect -12039 -4612 -11582 -4567
rect -12039 -4716 -11522 -4612
rect -7323 -4618 -6763 -4526
rect 6763 -4526 7400 -4497
rect 6763 -4618 7323 -4526
rect 11582 -4567 12095 -4464
rect 11582 -4612 12039 -4567
rect -7323 -4651 -6680 -4618
rect -11982 -4759 -11522 -4716
rect -7244 -4737 -6680 -4651
rect 6680 -4628 7323 -4618
rect 6680 -4737 9038 -4628
rect -11982 -4864 -11461 -4759
rect -7244 -4774 -6595 -4737
rect -11922 -4905 -11461 -4864
rect -7163 -4855 -6595 -4774
rect 6595 -4740 9038 -4737
rect 6595 -4774 7244 -4740
rect 6595 -4855 7163 -4774
rect -7163 -4897 -6508 -4855
rect -11922 -5012 -11397 -4905
rect -7080 -4939 -6508 -4897
rect -11861 -5050 -11397 -5012
rect -7266 -4971 -6508 -4939
rect 6508 -4897 7163 -4855
rect 6508 -4971 7080 -4897
rect -7266 -5029 -6419 -4971
rect -11861 -5159 -11332 -5050
rect -11797 -5195 -11332 -5159
rect -11797 -5305 -11265 -5195
rect -11732 -5339 -11265 -5305
rect -11732 -5450 -11197 -5339
rect -11665 -5481 -11197 -5450
rect -11665 -5595 -11126 -5481
rect -11597 -5623 -11126 -5595
rect -11597 -5739 -11054 -5623
rect -7266 -5638 -7176 -5029
rect -6995 -5086 -6419 -5029
rect 6419 -5018 7080 -4971
rect 6419 -5086 6995 -5018
rect 8926 -5046 9038 -4740
rect 11522 -4716 12039 -4612
rect 11522 -4759 11982 -4716
rect 11461 -4864 11982 -4759
rect 11461 -4905 11922 -4864
rect 11397 -5012 11922 -4905
rect 11397 -5050 11861 -5012
rect -6995 -5137 -6328 -5086
rect -6908 -5199 -6328 -5137
rect 6328 -5137 6995 -5086
rect 6328 -5199 6908 -5137
rect 11332 -5159 11861 -5050
rect 11332 -5172 11797 -5159
rect -6908 -5255 -6234 -5199
rect -6819 -5310 -6234 -5255
rect 6234 -5255 6908 -5199
rect 6234 -5310 6819 -5255
rect 10836 -5262 11797 -5172
rect -6819 -5371 -6139 -5310
rect -6728 -5420 -6139 -5371
rect 6139 -5371 6819 -5310
rect 11265 -5305 11797 -5262
rect 11265 -5339 11732 -5305
rect 6139 -5420 6728 -5371
rect -6728 -5486 -6042 -5420
rect -6634 -5528 -6042 -5486
rect 6042 -5486 6728 -5420
rect 11197 -5450 11732 -5339
rect 11197 -5481 11665 -5450
rect 11134 -5484 11665 -5481
rect 6042 -5528 6634 -5486
rect -6634 -5599 -5943 -5528
rect -11526 -5764 -11054 -5739
rect -8978 -5750 -7176 -5638
rect -6539 -5635 -5943 -5599
rect 5943 -5599 6634 -5528
rect 11126 -5595 11665 -5484
rect 5943 -5635 6539 -5599
rect 11126 -5623 11597 -5595
rect -6539 -5710 -5842 -5635
rect -11526 -5881 -10980 -5764
rect -11454 -5904 -10980 -5881
rect -11454 -6023 -10904 -5904
rect -11380 -6043 -10904 -6023
rect -11380 -6164 -10826 -6043
rect -8978 -6158 -8866 -5750
rect -7266 -5872 -7176 -5750
rect -6442 -5739 -5842 -5710
rect 5842 -5710 6539 -5635
rect 5842 -5739 6442 -5710
rect -6442 -5820 -5739 -5739
rect -6343 -5842 -5739 -5820
rect 5739 -5820 6442 -5739
rect 11054 -5739 11597 -5623
rect 11054 -5764 11526 -5739
rect 5739 -5842 6343 -5820
rect -6343 -5928 -5635 -5842
rect -6242 -5943 -5635 -5928
rect 5635 -5928 6343 -5842
rect 10980 -5881 11526 -5764
rect 10980 -5904 11454 -5881
rect 5635 -5943 6242 -5928
rect -6242 -6035 -5528 -5943
rect -6139 -6042 -5528 -6035
rect 5528 -6023 6242 -5943
rect 10904 -6023 11454 -5904
rect 5528 -6042 6930 -6023
rect -6139 -6139 -5420 -6042
rect 5420 -6113 6930 -6042
rect 10904 -6043 11380 -6023
rect 5420 -6139 6139 -6113
rect -11304 -6181 -10826 -6164
rect -11304 -6304 -10747 -6181
rect -9136 -6270 -8866 -6158
rect -6035 -6234 -5310 -6139
rect 5310 -6234 6035 -6139
rect -6035 -6242 -5199 -6234
rect -11226 -6318 -10747 -6304
rect -11226 -6443 -10666 -6318
rect -5928 -6328 -5199 -6242
rect 5199 -6242 6035 -6234
rect 5199 -6328 5928 -6242
rect -5928 -6343 -5086 -6328
rect -5820 -6419 -5086 -6343
rect 5086 -6343 5928 -6328
rect 5086 -6419 5820 -6343
rect -5820 -6442 -4971 -6419
rect -11147 -6455 -10666 -6443
rect -11147 -6581 -10583 -6455
rect -5710 -6508 -4971 -6442
rect 4971 -6442 5820 -6419
rect 4971 -6508 5710 -6442
rect -5710 -6539 -4855 -6508
rect -11066 -6589 -10583 -6581
rect -11066 -6718 -10499 -6589
rect -5599 -6595 -4855 -6539
rect 4855 -6539 5710 -6508
rect 4855 -6595 5599 -6539
rect -5599 -6634 -4737 -6595
rect -10983 -6723 -10499 -6718
rect -5486 -6680 -4737 -6634
rect 4737 -6634 5599 -6595
rect 4737 -6680 5486 -6634
rect -10983 -6855 -10413 -6723
rect -5486 -6728 -4618 -6680
rect -5371 -6763 -4618 -6728
rect 4618 -6728 5486 -6680
rect 4618 -6763 5371 -6728
rect -5371 -6819 -4497 -6763
rect -10899 -6856 -10413 -6855
rect -5255 -6844 -4497 -6819
rect 4497 -6819 5371 -6763
rect 4497 -6844 5255 -6819
rect -10899 -6988 -10325 -6856
rect -5255 -6908 -4374 -6844
rect -5137 -6923 -4374 -6908
rect 4374 -6908 5255 -6844
rect 4374 -6923 5137 -6908
rect -10899 -6989 -10235 -6988
rect -10813 -7119 -10235 -6989
rect -5137 -6995 -4251 -6923
rect -5018 -7000 -4251 -6995
rect 4251 -6995 5137 -6923
rect 6840 -6930 6930 -6113
rect 10826 -6164 11380 -6043
rect 10826 -6181 11304 -6164
rect 10747 -6304 11304 -6181
rect 10747 -6318 11226 -6304
rect 10666 -6443 11226 -6318
rect 10666 -6455 11147 -6443
rect 10583 -6581 11147 -6455
rect 10583 -6589 11066 -6581
rect 10499 -6718 11066 -6589
rect 10499 -6723 10983 -6718
rect 10413 -6855 10983 -6723
rect 10413 -6856 10899 -6855
rect 10325 -6988 10899 -6856
rect 10235 -6989 10899 -6988
rect 4251 -7000 5018 -6995
rect -5018 -7074 -4126 -7000
rect 4126 -7074 5018 -7000
rect -5018 -7080 -4000 -7074
rect -10813 -7123 -10144 -7119
rect -10725 -7248 -10144 -7123
rect -4897 -7146 -4000 -7080
rect 4000 -7080 5018 -7074
rect 4000 -7146 4897 -7080
rect 10235 -7119 10813 -6989
rect -4897 -7163 -3872 -7146
rect -4844 -7216 -3872 -7163
rect 3872 -7163 4897 -7146
rect 10144 -7123 10813 -7119
rect 3872 -7216 4774 -7163
rect -4844 -7244 -3743 -7216
rect -10725 -7256 -10051 -7248
rect -10635 -7376 -10051 -7256
rect -10635 -7388 -9957 -7376
rect -10544 -7503 -9957 -7388
rect -10544 -7519 -9861 -7503
rect -10451 -7629 -9861 -7519
rect -10451 -7648 -9763 -7629
rect -10357 -7754 -9763 -7648
rect -10357 -7776 -9664 -7754
rect -10261 -7877 -9664 -7776
rect -4844 -7806 -4754 -7244
rect -4651 -7284 -3743 -7244
rect 3743 -7244 4774 -7216
rect 3743 -7284 4651 -7244
rect 10144 -7248 10725 -7123
rect -4651 -7323 -3613 -7284
rect -4526 -7349 -3613 -7323
rect 3613 -7323 4651 -7284
rect 10051 -7256 10725 -7248
rect 3613 -7349 4526 -7323
rect -4526 -7400 -3482 -7349
rect -4400 -7412 -3482 -7400
rect 3482 -7400 4526 -7349
rect 10051 -7376 10635 -7256
rect 9957 -7388 10635 -7376
rect 3482 -7412 4400 -7400
rect -4400 -7473 -3349 -7412
rect 3349 -7473 4400 -7412
rect -4400 -7474 -3216 -7473
rect -4272 -7532 -3216 -7474
rect 3216 -7474 4400 -7473
rect 3216 -7532 4272 -7474
rect 9957 -7503 10544 -7388
rect -4272 -7546 -3082 -7532
rect -4143 -7588 -3082 -7546
rect 3082 -7546 4272 -7532
rect 9861 -7519 10544 -7503
rect 3082 -7588 4187 -7546
rect -4143 -7616 -2946 -7588
rect -4013 -7642 -2946 -7616
rect 2946 -7616 4187 -7588
rect 2946 -7642 4013 -7616
rect -4013 -7684 -2810 -7642
rect -3882 -7693 -2810 -7684
rect 2810 -7684 4013 -7642
rect 2810 -7693 3882 -7684
rect -3882 -7742 -2672 -7693
rect 2672 -7742 3882 -7693
rect -3882 -7749 -2534 -7742
rect -3749 -7788 -2534 -7749
rect 2534 -7749 3882 -7742
rect 4097 -7689 4187 -7616
rect 9861 -7629 10451 -7519
rect 9763 -7648 10451 -7629
rect 2534 -7788 3749 -7749
rect 4097 -7779 4244 -7689
rect 9763 -7754 10357 -7648
rect 9664 -7756 10357 -7754
rect -3749 -7812 -2395 -7788
rect -3616 -7832 -2395 -7812
rect 2395 -7812 3749 -7788
rect 2395 -7832 3616 -7812
rect -3616 -7873 -2255 -7832
rect -3482 -7874 -2255 -7873
rect 2255 -7873 3616 -7832
rect 2255 -7874 3482 -7873
rect -10261 -7903 -9563 -7877
rect -10163 -7999 -9563 -7903
rect -3482 -7913 -2115 -7874
rect 2115 -7913 3482 -7874
rect -3482 -7932 -1974 -7913
rect -3346 -7950 -1974 -7932
rect 1974 -7932 3482 -7913
rect 1974 -7950 3346 -7932
rect -3346 -7984 -1832 -7950
rect 1832 -7984 3346 -7950
rect -3346 -7988 -1689 -7984
rect -10163 -8029 -9461 -7999
rect -10064 -8120 -9461 -8029
rect -3210 -8016 -1689 -7988
rect 1689 -7988 3346 -7984
rect 1689 -8016 3210 -7988
rect -3210 -8042 -1546 -8016
rect -3072 -8045 -1546 -8042
rect 1546 -8042 3210 -8016
rect 1546 -8045 3072 -8042
rect -3072 -8072 -1402 -8045
rect 1402 -8072 3072 -8045
rect -3072 -8093 -1258 -8072
rect -2934 -8096 -1258 -8093
rect 1258 -8093 3072 -8072
rect 1258 -8096 2934 -8093
rect -2934 -8118 -1114 -8096
rect 1114 -8118 2934 -8096
rect -10064 -8154 -9357 -8120
rect -2934 -8137 -969 -8118
rect 969 -8137 2934 -8118
rect -2934 -8142 -823 -8137
rect -9963 -8239 -9357 -8154
rect -2795 -8153 -823 -8142
rect 823 -8142 2934 -8137
rect 823 -8153 2795 -8142
rect -2795 -8168 -678 -8153
rect 678 -8168 2795 -8153
rect -2795 -8179 -532 -8168
rect 532 -8179 2795 -8168
rect -2795 -8188 -385 -8179
rect 385 -8188 2795 -8179
rect -2655 -8194 -239 -8188
rect 239 -8194 2655 -8188
rect -2655 -8198 -93 -8194
rect 93 -8198 2655 -8194
rect -2655 -8232 2655 -8198
rect -9963 -8277 -9252 -8239
rect -2515 -8274 2515 -8232
rect -9861 -8357 -9252 -8277
rect -2374 -8313 2374 -8274
rect -2232 -8350 2232 -8313
rect -9861 -8399 -9145 -8357
rect -2089 -8384 2089 -8350
rect -9757 -8474 -9145 -8399
rect -1958 -8416 1946 -8384
rect -9757 -8520 -9037 -8474
rect -9652 -8589 -9037 -8520
rect -9652 -8639 -8927 -8589
rect -9545 -8703 -8927 -8639
rect -9545 -8757 -8816 -8703
rect -9437 -8816 -8816 -8757
rect -9437 -8874 -8703 -8816
rect -9327 -8927 -8703 -8874
rect -9327 -8989 -8589 -8927
rect -9216 -9037 -8589 -8989
rect -9216 -9103 -8474 -9037
rect -9103 -9145 -8474 -9103
rect -9103 -9216 -8357 -9145
rect -8989 -9252 -8357 -9216
rect -8989 -9327 -8239 -9252
rect -8874 -9357 -8239 -9327
rect -8874 -9437 -8120 -9357
rect -8757 -9461 -8120 -9437
rect -8757 -9545 -7999 -9461
rect -8639 -9563 -7999 -9545
rect -8639 -9652 -7877 -9563
rect -8520 -9664 -7877 -9652
rect -8520 -9757 -7754 -9664
rect -8399 -9763 -7754 -9757
rect -8399 -9861 -7629 -9763
rect -8277 -9957 -7503 -9861
rect -8277 -9963 -7376 -9957
rect -8154 -10051 -7376 -9963
rect -7266 -10051 -7176 -8672
rect -1958 -8938 -1868 -8416
rect -1802 -8445 1802 -8416
rect -1658 -8472 1658 -8445
rect -1514 -8496 1514 -8472
rect -1369 -8518 1369 -8496
rect -1223 -8537 1223 -8518
rect -1078 -8553 1078 -8537
rect -932 -8568 932 -8553
rect -785 -8579 785 -8568
rect -639 -8588 639 -8579
rect -493 -8594 493 -8588
rect -346 -8598 346 -8594
rect -200 -8600 199 -8598
rect 1132 -9170 1222 -8537
rect 4154 -8581 4244 -7779
rect 8948 -7776 10357 -7756
rect 8948 -7846 10261 -7776
rect 9664 -7877 10261 -7846
rect 9563 -7903 10261 -7877
rect 9563 -7999 10163 -7903
rect 9461 -8029 10163 -7999
rect 9461 -8120 10064 -8029
rect 9357 -8154 10064 -8120
rect 9357 -8239 9963 -8154
rect 9252 -8277 9963 -8239
rect 9252 -8357 9861 -8277
rect 9145 -8399 9861 -8357
rect 9145 -8474 9757 -8399
rect 9037 -8520 9757 -8474
rect 9037 -8589 9652 -8520
rect 8927 -8639 9652 -8589
rect 8927 -8703 9545 -8639
rect 8816 -8757 9545 -8703
rect 8816 -8816 9437 -8757
rect 8703 -8874 9437 -8816
rect 8703 -8927 9327 -8874
rect 8589 -8989 9327 -8927
rect 8589 -9037 9216 -8989
rect 8474 -9103 9216 -9037
rect 8474 -9145 9103 -9103
rect 8357 -9216 9103 -9145
rect 8357 -9252 8989 -9216
rect 8239 -9327 8989 -9252
rect 8239 -9357 8874 -9327
rect 8120 -9437 8874 -9357
rect 8120 -9461 8757 -9437
rect 7999 -9545 8757 -9461
rect 7999 -9563 8639 -9545
rect 7877 -9652 8639 -9563
rect 7877 -9664 8520 -9652
rect -8154 -10064 -7176 -10051
rect -8029 -10144 -7176 -10064
rect -8029 -10163 -7119 -10144
rect -7903 -10235 -7119 -10163
rect -7903 -10261 -6988 -10235
rect -7776 -10325 -6988 -10261
rect 6840 -10325 6930 -9730
rect 7754 -9757 8520 -9664
rect 7754 -9763 8399 -9757
rect 7629 -9861 8399 -9763
rect 7503 -9957 8277 -9861
rect 7376 -9963 8277 -9957
rect 7376 -10051 8154 -9963
rect 7248 -10064 8154 -10051
rect 7248 -10144 8029 -10064
rect 7119 -10163 8029 -10144
rect 7119 -10235 7903 -10163
rect 6988 -10261 7903 -10235
rect 6988 -10325 7776 -10261
rect -7776 -10357 -6856 -10325
rect -7648 -10413 -6856 -10357
rect 6840 -10357 7776 -10325
rect 6840 -10413 7648 -10357
rect -7648 -10451 -6723 -10413
rect -7519 -10499 -6723 -10451
rect 6723 -10451 7648 -10413
rect 6723 -10499 7519 -10451
rect -7519 -10544 -6589 -10499
rect -7388 -10583 -6589 -10544
rect 6589 -10544 7519 -10499
rect 6589 -10583 7388 -10544
rect -7388 -10635 -6455 -10583
rect -7256 -10666 -6455 -10635
rect -7256 -10725 -6318 -10666
rect -7123 -10747 -6318 -10725
rect -7123 -10813 -6181 -10747
rect -6989 -10826 -6181 -10813
rect -6989 -10899 -6043 -10826
rect -6855 -10904 -6043 -10899
rect -6855 -10980 -5904 -10904
rect -6855 -10983 -5764 -10980
rect -6718 -11054 -5764 -10983
rect -6718 -11066 -5623 -11054
rect -6581 -11126 -5623 -11066
rect -6581 -11147 -5481 -11126
rect -6443 -11197 -5481 -11147
rect -6443 -11226 -5339 -11197
rect -6304 -11265 -5339 -11226
rect -6304 -11304 -5195 -11265
rect -6164 -11332 -5195 -11304
rect -6164 -11380 -5050 -11332
rect -6023 -11397 -5050 -11380
rect -6023 -11454 -4905 -11397
rect -5881 -11461 -4905 -11454
rect -4844 -11461 -4754 -10606
rect 6455 -10635 7388 -10583
rect 6455 -10666 7256 -10635
rect 6318 -10725 7256 -10666
rect 6318 -10747 7123 -10725
rect 6181 -10813 7123 -10747
rect 6181 -10826 6989 -10813
rect 6043 -10899 6989 -10826
rect 6043 -10904 6855 -10899
rect 5904 -10980 6855 -10904
rect 5764 -10983 6855 -10980
rect 5764 -11054 6718 -10983
rect 5623 -11066 6718 -11054
rect 5623 -11126 6581 -11066
rect 5481 -11147 6581 -11126
rect -5881 -11522 -4754 -11461
rect -5881 -11526 -4612 -11522
rect -5739 -11582 -4612 -11526
rect -5739 -11597 -4464 -11582
rect -5595 -11639 -4464 -11597
rect -5595 -11665 -4316 -11639
rect -5450 -11695 -4316 -11665
rect 4154 -11695 4244 -11173
rect 5481 -11197 6443 -11147
rect 5339 -11226 6443 -11197
rect 5339 -11265 6304 -11226
rect 5195 -11304 6304 -11265
rect 5195 -11332 6164 -11304
rect 5050 -11380 6164 -11332
rect 5050 -11397 6023 -11380
rect 4905 -11454 6023 -11397
rect 4905 -11461 5881 -11454
rect 4759 -11522 5881 -11461
rect 4612 -11526 5881 -11522
rect 4612 -11582 5739 -11526
rect 4464 -11597 5739 -11582
rect 4464 -11639 5595 -11597
rect 4316 -11665 5595 -11639
rect 4316 -11695 5450 -11665
rect -5450 -11732 -4167 -11695
rect -5305 -11749 -4167 -11732
rect 4154 -11732 5450 -11695
rect -5305 -11797 -4017 -11749
rect -5159 -11801 -4017 -11797
rect -5159 -11851 -3866 -11801
rect -5159 -11861 -3715 -11851
rect -5012 -11900 -3715 -11861
rect -5012 -11922 -3564 -11900
rect -4864 -11946 -3564 -11922
rect -4864 -11982 -3411 -11946
rect -4716 -11990 -3411 -11982
rect -4716 -12033 -3258 -11990
rect -4716 -12039 -3105 -12033
rect -4567 -12073 -3105 -12039
rect -4567 -12095 -2951 -12073
rect -4417 -12112 -2951 -12095
rect -4417 -12149 -2796 -12112
rect -4266 -12183 -2641 -12149
rect -4266 -12201 -2486 -12183
rect -4115 -12216 -2486 -12201
rect -4115 -12247 -2330 -12216
rect -4115 -12251 -2174 -12247
rect -3964 -12276 -2174 -12251
rect -3964 -12300 -2017 -12276
rect -3811 -12303 -2017 -12300
rect -1958 -12303 -1868 -11738
rect 4154 -11749 5305 -11732
rect 4017 -11797 5305 -11749
rect 4017 -11801 5159 -11797
rect 3866 -11851 5159 -11801
rect 3715 -11861 5159 -11851
rect 3715 -11900 5012 -11861
rect 3564 -11922 5012 -11900
rect 3564 -11946 4864 -11922
rect -3811 -12328 -1860 -12303
rect 1132 -12309 1222 -11970
rect 3411 -11982 4864 -11946
rect 3411 -11990 4716 -11982
rect 3258 -12033 4716 -11990
rect 3105 -12039 4716 -12033
rect 3105 -12073 4567 -12039
rect 2951 -12095 4567 -12073
rect 2951 -12112 4417 -12095
rect 2796 -12149 4417 -12112
rect 2641 -12183 4266 -12149
rect 2486 -12201 4266 -12183
rect 2486 -12216 4115 -12201
rect 2330 -12247 4115 -12216
rect 2174 -12251 4115 -12247
rect 2174 -12276 3964 -12251
rect 2017 -12300 3964 -12276
rect 2017 -12303 3811 -12300
rect -3811 -12346 -1703 -12328
rect -3658 -12351 -1703 -12346
rect -3658 -12372 -1546 -12351
rect -3658 -12390 -1388 -12372
rect -3505 -12391 -1388 -12390
rect 1132 -12391 1277 -12309
rect 1860 -12328 3811 -12303
rect 1703 -12346 3811 -12328
rect 1703 -12351 3658 -12346
rect 1546 -12372 3658 -12351
rect 1388 -12390 3658 -12372
rect 1388 -12391 3505 -12390
rect -3505 -12408 -1230 -12391
rect 1132 -12408 3505 -12391
rect -3505 -12423 -1071 -12408
rect 1071 -12423 3505 -12408
rect -3505 -12433 -913 -12423
rect -3351 -12435 -913 -12433
rect 913 -12433 3505 -12423
rect 913 -12435 3351 -12433
rect -3351 -12446 -754 -12435
rect 754 -12446 3351 -12435
rect -3351 -12455 -595 -12446
rect 595 -12455 3351 -12446
rect -3351 -12462 -436 -12455
rect 436 -12462 3351 -12455
rect -3351 -12467 -277 -12462
rect 277 -12467 3351 -12462
rect -3351 -12470 -118 -12467
rect 118 -12470 3351 -12467
rect -3351 -12473 3351 -12470
rect -3196 -12512 3196 -12473
rect -3041 -12549 3041 -12512
rect -2886 -12583 2886 -12549
rect -2730 -12616 2730 -12583
rect -2574 -12647 2574 -12616
rect -2417 -12676 2417 -12647
rect -2260 -12703 2260 -12676
rect -2103 -12728 2103 -12703
rect -1946 -12751 1946 -12728
rect -1788 -12772 1788 -12751
rect -1630 -12791 1630 -12772
rect -1471 -12808 1471 -12791
rect -1313 -12823 1313 -12808
rect -1154 -12835 1154 -12823
rect -995 -12846 995 -12835
rect -836 -12855 836 -12846
rect -677 -12862 677 -12855
rect -518 -12867 518 -12862
rect -359 -12870 359 -12867
rect -200 -12872 199 -12870
use skullfet_inverter_5v  skullfet_inverter_0
timestamp 1735290363
transform 1 0 9800 0 1 -2000
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_1
timestamp 1735290363
transform -1 0 11536 0 1 1384
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_2
timestamp 1735290363
transform 1 0 7592 0 1 4458
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_3
timestamp 1735290363
transform 1 0 5484 0 1 6730
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_4
timestamp 1735290363
transform 1 0 2798 0 1 8280
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_5
timestamp 1735290363
transform 1 0 -224 0 1 8970
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_6
timestamp 1735290363
transform 1 0 -3314 0 1 8738
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_7
timestamp 1735290363
transform 1 0 -6198 0 1 7606
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_8
timestamp 1735290363
transform 1 0 -8622 0 1 5672
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_9
timestamp 1735290363
transform 1 0 -10370 0 1 3512
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_10
timestamp 1735290363
transform 1 0 -11282 0 1 150
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_11
timestamp 1735290363
transform 1 0 -12082 0 1 -3150
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_12
timestamp 1735290363
transform -1 0 -8470 0 1 -6512
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_13
timestamp 1735290363
transform -1 0 -6622 0 -1 -5672
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_14
timestamp 1735290363
transform -1 0 -4200 0 -1 -7606
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_15
timestamp 1735290363
transform -1 0 -1314 0 -1 -8738
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_16
timestamp 1735290363
transform -1 0 1776 0 -1 -8970
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_17
timestamp 1735290363
transform -1 0 4798 0 -1 -8280
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_18
timestamp 1735290363
transform -1 0 7484 0 -1 -6730
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_19
timestamp 1735290363
transform -1 0 9592 0 -1 -4758
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_20
timestamp 1735290363
transform -1 0 11480 0 -1 -2174
box 454 132 2110 3088
<< end >>
