magic
tech sky130A
magscale 1 2
timestamp 1735333972
<< metal1 >>
rect 18107 44173 18354 44269
rect 18450 44173 18460 44269
rect 12286 43628 12304 43724
rect 12400 43628 12652 43724
rect 13432 43226 13442 43338
rect 13554 43226 13564 43338
rect 12010 43089 12020 43145
rect 12130 43089 12140 43145
rect 10430 42937 10440 43037
rect 10540 42937 10550 43037
rect 12024 34460 12124 41646
rect 1494 22582 1504 22882
rect 1804 22582 1814 22882
rect 6142 22866 6152 23106
rect 6352 22866 6362 23106
<< via1 >>
rect 18354 44173 18450 44269
rect 12304 43628 12400 43724
rect 13442 43226 13554 43338
rect 12020 43089 12130 43145
rect 10440 42937 10540 43037
rect 1504 22582 1804 22882
rect 6152 22866 6352 23106
<< metal2 >>
rect 17172 44818 17236 44828
rect 17172 44728 17236 44738
rect 17724 44818 17788 44828
rect 17724 44728 17788 44738
rect 18276 44818 18340 44828
rect 17174 44554 17226 44728
rect 12866 44502 17226 44554
rect 12866 43760 12918 44502
rect 17728 44450 17780 44728
rect 14808 44398 17780 44450
rect 14808 43752 14860 44398
rect 18276 44366 18340 44738
rect 16736 44314 18340 44366
rect 16736 43772 16788 44314
rect 18354 44269 18450 44279
rect 18354 44163 18450 44173
rect 18080 43980 18140 43990
rect 18080 43890 18140 43900
rect 12282 43724 12420 43746
rect 12282 43628 12304 43724
rect 12400 43628 12420 43724
rect 12282 43606 12420 43628
rect 13442 43338 13554 43348
rect 12020 43145 12130 43155
rect 12020 43079 12130 43089
rect 10440 43037 10540 43047
rect 10540 42937 10732 43026
rect 10440 42936 10732 42937
rect 10440 42927 10540 42936
rect 13442 42914 13554 43226
rect 6152 23106 6352 23116
rect 1504 22882 1804 22892
rect 6152 22856 6352 22866
rect 1504 22572 1804 22582
<< via2 >>
rect 17172 44738 17236 44818
rect 17724 44738 17788 44818
rect 18276 44738 18340 44818
rect 18354 44173 18450 44269
rect 18080 43900 18140 43980
rect 12304 43628 12400 43724
rect 13442 43226 13554 43338
rect 12020 43089 12130 43145
rect 10440 42937 10540 43037
rect 1504 22582 1804 22882
rect 6152 22866 6352 23106
<< metal3 >>
rect 17162 44818 17246 44853
rect 17162 44738 17172 44818
rect 17236 44738 17246 44818
rect 17162 44733 17246 44738
rect 17714 44818 17798 44853
rect 17714 44738 17724 44818
rect 17788 44738 17798 44818
rect 17714 44733 17798 44738
rect 18266 44818 18350 44853
rect 18266 44738 18276 44818
rect 18340 44738 18350 44818
rect 18266 44733 18350 44738
rect 18344 44272 18460 44274
rect 18312 44269 18512 44272
rect 18312 44173 18354 44269
rect 18450 44173 18512 44269
rect 18060 43980 18160 44000
rect 18060 43900 18078 43980
rect 18142 43900 18160 43980
rect 18060 43880 18160 43900
rect 12282 43729 12420 43746
rect 12282 43623 12299 43729
rect 12405 43623 12420 43729
rect 12282 43606 12420 43623
rect 18312 43410 18512 44173
rect 624 43408 18512 43410
rect 624 43210 658 43408
rect 648 43208 658 43210
rect 858 43338 18512 43408
rect 858 43226 13442 43338
rect 13554 43226 18512 43338
rect 858 43210 18512 43226
rect 858 43208 868 43210
rect 11986 43086 11996 43150
rect 12146 43086 12156 43150
rect 12010 43084 12140 43086
rect 10430 43037 10550 43042
rect 10430 42937 10440 43037
rect 10540 42937 10550 43037
rect 10430 42932 10550 42937
rect 6142 23106 6362 23111
rect 106 22466 116 22974
rect 524 22882 554 22974
rect 1494 22882 1814 22887
rect 524 22582 1504 22882
rect 1804 22582 1814 22882
rect 6142 22866 6152 23106
rect 6352 22866 6362 23106
rect 6142 22861 6362 22866
rect 524 22466 554 22582
rect 1494 22577 1814 22582
<< via3 >>
rect 17172 44738 17236 44818
rect 17724 44738 17788 44818
rect 18276 44738 18340 44818
rect 18078 43900 18080 43980
rect 18080 43900 18140 43980
rect 18140 43900 18142 43980
rect 12299 43724 12405 43729
rect 12299 43628 12304 43724
rect 12304 43628 12400 43724
rect 12400 43628 12405 43724
rect 12299 43623 12405 43628
rect 658 43208 858 43408
rect 11996 43145 12146 43150
rect 11996 43089 12020 43145
rect 12020 43089 12130 43145
rect 12130 43089 12146 43145
rect 11996 43086 12146 43089
rect 10440 42937 10540 43037
rect 116 22466 524 22974
rect 6152 22866 6352 23106
<< metal4 >>
rect 6134 44610 6194 45152
rect 6686 44610 6746 45152
rect 7238 44610 7298 45152
rect 7790 44610 7850 45152
rect 8342 44610 8402 45152
rect 8894 44610 8954 45152
rect 9446 44610 9506 45152
rect 9998 44610 10058 45152
rect 10550 44610 10610 45152
rect 11102 44610 11162 45152
rect 11654 44610 11714 45152
rect 12206 44610 12266 45152
rect 12758 44610 12818 45152
rect 13310 44610 13370 45152
rect 13862 44610 13922 45152
rect 14414 44610 14474 45152
rect 14966 44610 15026 45152
rect 15518 44610 15578 45152
rect 16070 44610 16130 45152
rect 16622 44610 16682 45152
rect 17174 44819 17234 45152
rect 17726 44819 17786 45152
rect 18278 44819 18338 45152
rect 17171 44818 17237 44819
rect 17171 44738 17172 44818
rect 17236 44738 17237 44818
rect 17171 44737 17237 44738
rect 17723 44818 17789 44819
rect 17723 44738 17724 44818
rect 17788 44738 17789 44818
rect 17723 44737 17789 44738
rect 18275 44818 18341 44819
rect 18275 44738 18276 44818
rect 18340 44738 18341 44818
rect 18275 44737 18341 44738
rect 200 44410 16682 44610
rect 18830 44422 18890 45152
rect 19382 44952 19442 45152
rect 19934 44952 19994 45152
rect 20486 44952 20546 45152
rect 21038 44952 21098 45152
rect 21590 44952 21650 45152
rect 22142 44952 22202 45152
rect 22694 44952 22754 45152
rect 23246 44952 23306 45152
rect 23798 44952 23858 45152
rect 24350 44952 24410 45152
rect 24902 44952 24962 45152
rect 25454 44952 25514 45152
rect 26006 44952 26066 45152
rect 26558 44952 26618 45152
rect 27110 44952 27170 45152
rect 27662 44952 27722 45152
rect 28214 44952 28274 45152
rect 28766 44952 28826 45152
rect 29318 44952 29378 45152
rect 200 22975 500 44410
rect 600 43408 900 44152
rect 600 43208 658 43408
rect 858 43208 900 43408
rect 115 22974 538 22975
rect 115 22466 116 22974
rect 524 22466 538 22974
rect 115 22465 538 22466
rect 200 1000 500 22465
rect 600 1000 900 43208
rect 1000 23122 1300 44152
rect 10475 43038 10545 44410
rect 12098 43730 12298 44410
rect 18082 44362 18890 44422
rect 18082 44000 18142 44362
rect 18060 43980 18160 44000
rect 18060 43900 18078 43980
rect 18142 43900 18160 43980
rect 18060 43880 18160 43900
rect 12098 43729 12406 43730
rect 12098 43628 12299 43729
rect 12298 43623 12299 43628
rect 12405 43623 12406 43729
rect 12298 43622 12406 43623
rect 18082 43514 18142 43880
rect 12034 43454 18142 43514
rect 12034 43151 12094 43454
rect 11995 43150 12147 43151
rect 11995 43086 11996 43150
rect 12146 43086 12147 43150
rect 11995 43085 12147 43086
rect 10439 43037 10545 43038
rect 10439 42937 10440 43037
rect 10540 42937 10545 43037
rect 10439 42936 10541 42937
rect 1000 23106 6384 23122
rect 1000 22866 6152 23106
rect 6352 22866 6384 23106
rect 1000 22822 6384 22866
rect 1000 1000 1300 22822
rect 27234 0 27414 200 0
rect 23370 0 23550 200 0
rect 19506 0 19686 200 0
rect 15642 0 15822 200 0
rect 11778 0 11958 200 0
rect 7914 0 8094 200 0
rect 4050 0 4230 200 0
rect 186 0 366 200 0
use big_skull  big_skull_0
timestamp 1713168785
transform 1 0 9474 0 1 33040
box 1040 -17680 11960 -2080
use freq_divider  freq_divider_0
timestamp 1725542573
transform -1 0 22072 0 1 43628
box 3864 0 9552 640
use ring  ring_0
timestamp 1735296899
transform 1 0 16088 0 1 22922
box -14600 -14600 14600 14600
use skullfet_inverter_5v  skullfet_level_shifter
timestamp 1735290363
transform 0 -1 13730 -1 0 43580
box 454 132 2110 3088
<< labels >>
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 240 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 29318 44952 29378 45152 0 FreeSans 240 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 28214 44952 28274 45152 0 FreeSans 240 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27662 44952 27722 45152 0 FreeSans 240 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 27110 44952 27170 45152 0 FreeSans 240 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 240 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 26006 44952 26066 45152 0 FreeSans 240 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 25454 44952 25514 45152 0 FreeSans 240 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 24902 44952 24962 45152 0 FreeSans 240 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 240 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 23798 44952 23858 45152 0 FreeSans 240 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 23246 44952 23306 45152 0 FreeSans 240 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 22694 44952 22754 45152 0 FreeSans 240 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 240 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 21590 44952 21650 45152 0 FreeSans 240 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 21038 44952 21098 45152 0 FreeSans 240 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 20486 44952 20546 45152 0 FreeSans 240 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 240 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19382 44952 19442 45152 0 FreeSans 240 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 9998 44952 10058 45152 0 FreeSans 240 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 9446 44952 9506 45152 0 FreeSans 240 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 240 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 8342 44952 8402 45152 0 FreeSans 240 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 7790 44952 7850 45152 0 FreeSans 240 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 7238 44952 7298 45152 0 FreeSans 240 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 240 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 6134 44952 6194 45152 0 FreeSans 240 90 0 0 uio_oe[7]
port 26 nsew signal output
flabel metal4 s 14414 44952 14474 45152 0 FreeSans 240 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 13862 44952 13922 45152 0 FreeSans 240 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 240 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 12758 44952 12818 45152 0 FreeSans 240 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 12206 44952 12266 45152 0 FreeSans 240 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 11654 44952 11714 45152 0 FreeSans 240 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 240 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 10550 44952 10610 45152 0 FreeSans 240 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 18830 44952 18890 45152 0 FreeSans 240 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 18278 44952 18338 45152 0 FreeSans 240 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 240 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 17174 44952 17234 45152 0 FreeSans 240 90 0 0 uo_out[3]
port 38 nsew signal output
flabel metal4 s 16622 44952 16682 45152 0 FreeSans 240 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 16070 44952 16130 45152 0 FreeSans 240 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 240 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 14966 44952 15026 45152 0 FreeSans 240 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 43 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 44 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 45 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 46 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 47 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 48 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 49 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 50 nsew signal bidirectional
flabel metal4 1000 1000 1300 44152 1 FreeSans 2 0 0 0 VAPWR
port 51 nsew power bidirectional
flabel metal4 600 1000 900 44152 1 FreeSans 2 0 0 0 VDPWR
port 52 nsew power bidirectional
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VGND
port 53 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
