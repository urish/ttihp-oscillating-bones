magic
tech sky130A
timestamp 1713168785
<< metal4 >>
rect 1989 -1105 3757 -884
rect 1768 -1326 3757 -1105
rect 1326 -1768 4199 -1326
rect 1105 -2652 4420 -1768
rect 1105 -2873 1768 -2652
rect 3757 -2873 4420 -2652
rect 2431 -3315 3094 -2652
rect 1105 -3094 1547 -2873
rect 3978 -3094 4420 -2873
rect 1326 -3757 1547 -3094
rect 2210 -3536 3315 -3315
rect 3978 -3536 4199 -3094
rect 1547 -3757 1768 -3315
rect 1989 -4420 2431 -3536
rect 1768 -3978 1989 -3536
rect 2431 -3757 2652 -3536
rect 3757 -3978 3978 -3315
rect 2873 -3757 3757 -3536
rect 3094 -3978 3757 -3757
rect 2431 -4420 3536 -3978
rect 1989 -4641 2210 -4420
rect 2431 -4641 2652 -4420
rect 2873 -4641 3094 -4420
rect 3315 -4641 3536 -4420
rect 663 -7514 884 -7293
rect 442 -7293 1105 -7072
rect 442 -7072 1326 -6851
rect 442 -6851 1768 -6630
rect 663 -6630 2210 -6409
rect 1768 -6409 2652 -6188
rect 2873 -6409 3757 -6188
rect 3315 -6630 5083 -6409
rect 3757 -6851 5083 -6630
rect 4199 -7072 5083 -6851
rect 4420 -7293 5083 -7072
rect 4641 -7514 4862 -7293
rect 2210 -6188 3315 -5746
rect 1768 -5746 2652 -5525
rect 2873 -5746 3757 -5525
rect 1326 -5525 2210 -5304
rect 3315 -5525 4199 -5304
rect 663 -5304 1989 -5083
rect 3536 -5304 4862 -5083
rect 442 -5083 1547 -4641
rect 3978 -5083 5083 -4641
rect 663 -4641 1326 -4420
rect 4199 -4641 4862 -4420
<< metal3 >>
rect 1989 -1105 3757 -884
rect 1768 -1326 3757 -1105
rect 1326 -1768 4199 -1326
rect 1105 -2652 4420 -1768
rect 1105 -2873 1768 -2652
rect 3757 -2873 4420 -2652
rect 2431 -3315 3094 -2652
rect 1105 -3094 1547 -2873
rect 3978 -3094 4420 -2873
rect 1326 -3757 1547 -3094
rect 2210 -3536 3315 -3315
rect 3978 -3536 4199 -3094
rect 1547 -3757 1768 -3315
rect 1989 -4420 2431 -3536
rect 1768 -3978 1989 -3536
rect 2431 -3757 2652 -3536
rect 3757 -3978 3978 -3315
rect 2873 -3757 3757 -3536
rect 3094 -3978 3757 -3757
rect 2431 -4420 3536 -3978
rect 1989 -4641 2210 -4420
rect 2431 -4641 2652 -4420
rect 2873 -4641 3094 -4420
rect 3315 -4641 3536 -4420
rect 663 -7514 884 -7293
rect 442 -7293 1105 -7072
rect 442 -7072 1326 -6851
rect 442 -6851 1768 -6630
rect 663 -6630 2210 -6409
rect 1768 -6409 2652 -6188
rect 2873 -6409 3757 -6188
rect 3315 -6630 5083 -6409
rect 3757 -6851 5083 -6630
rect 4199 -7072 5083 -6851
rect 4420 -7293 5083 -7072
rect 4641 -7514 4862 -7293
rect 2210 -6188 3315 -5746
rect 1768 -5746 2652 -5525
rect 2873 -5746 3757 -5525
rect 1326 -5525 2210 -5304
rect 3315 -5525 4199 -5304
rect 663 -5304 1989 -5083
rect 3536 -5304 4862 -5083
rect 442 -5083 1547 -4641
rect 3978 -5083 5083 -4641
rect 663 -4641 1326 -4420
rect 4199 -4641 4862 -4420
<< metal2 >>
rect 1989 -1105 3757 -884
rect 1768 -1326 3757 -1105
rect 1326 -1768 4199 -1326
rect 1105 -2652 4420 -1768
rect 1105 -2873 1768 -2652
rect 3757 -2873 4420 -2652
rect 2431 -3315 3094 -2652
rect 1105 -3094 1547 -2873
rect 3978 -3094 4420 -2873
rect 1326 -3757 1547 -3094
rect 2210 -3536 3315 -3315
rect 3978 -3536 4199 -3094
rect 1547 -3757 1768 -3315
rect 1989 -4420 2431 -3536
rect 1768 -3978 1989 -3536
rect 2431 -3757 2652 -3536
rect 3757 -3978 3978 -3315
rect 2873 -3757 3757 -3536
rect 3094 -3978 3757 -3757
rect 2431 -4420 3536 -3978
rect 1989 -4641 2210 -4420
rect 2431 -4641 2652 -4420
rect 2873 -4641 3094 -4420
rect 3315 -4641 3536 -4420
rect 663 -7514 884 -7293
rect 442 -7293 1105 -7072
rect 442 -7072 1326 -6851
rect 442 -6851 1768 -6630
rect 663 -6630 2210 -6409
rect 1768 -6409 2652 -6188
rect 2873 -6409 3757 -6188
rect 3315 -6630 5083 -6409
rect 3757 -6851 5083 -6630
rect 4199 -7072 5083 -6851
rect 4420 -7293 5083 -7072
rect 4641 -7514 4862 -7293
rect 2210 -6188 3315 -5746
rect 1768 -5746 2652 -5525
rect 2873 -5746 3757 -5525
rect 1326 -5525 2210 -5304
rect 3315 -5525 4199 -5304
rect 663 -5304 1989 -5083
rect 3536 -5304 4862 -5083
rect 442 -5083 1547 -4641
rect 3978 -5083 5083 -4641
rect 663 -4641 1326 -4420
rect 4199 -4641 4862 -4420
<< metal1 >>
rect 1989 -1105 3757 -884
rect 1768 -1326 3757 -1105
rect 1326 -1768 4199 -1326
rect 1105 -2652 4420 -1768
rect 1105 -2873 1768 -2652
rect 3757 -2873 4420 -2652
rect 2431 -3315 3094 -2652
rect 1105 -3094 1547 -2873
rect 3978 -3094 4420 -2873
rect 1326 -3757 1547 -3094
rect 2210 -3536 3315 -3315
rect 3978 -3536 4199 -3094
rect 1547 -3757 1768 -3315
rect 1989 -4420 2431 -3536
rect 1768 -3978 1989 -3536
rect 2431 -3757 2652 -3536
rect 3757 -3978 3978 -3315
rect 2873 -3757 3757 -3536
rect 3094 -3978 3757 -3757
rect 2431 -4420 3536 -3978
rect 1989 -4641 2210 -4420
rect 2431 -4641 2652 -4420
rect 2873 -4641 3094 -4420
rect 3315 -4641 3536 -4420
rect 663 -7514 884 -7293
rect 442 -7293 1105 -7072
rect 442 -7072 1326 -6851
rect 442 -6851 1768 -6630
rect 663 -6630 2210 -6409
rect 1768 -6409 2652 -6188
rect 2873 -6409 3757 -6188
rect 3315 -6630 5083 -6409
rect 3757 -6851 5083 -6630
rect 4199 -7072 5083 -6851
rect 4420 -7293 5083 -7072
rect 4641 -7514 4862 -7293
rect 2210 -6188 3315 -5746
rect 1768 -5746 2652 -5525
rect 2873 -5746 3757 -5525
rect 1326 -5525 2210 -5304
rect 3315 -5525 4199 -5304
rect 663 -5304 1989 -5083
rect 3536 -5304 4862 -5083
rect 442 -5083 1547 -4641
rect 3978 -5083 5083 -4641
rect 663 -4641 1326 -4420
rect 4199 -4641 4862 -4420
<< fillblock >>
rect 1989 -1105 3757 -884
rect 1768 -1326 3757 -1105
rect 1326 -1768 4199 -1326
rect 1105 -2652 4420 -1768
rect 1105 -2873 1768 -2652
rect 3757 -2873 4420 -2652
rect 2431 -3315 3094 -2652
rect 1105 -3094 1547 -2873
rect 3978 -3094 4420 -2873
rect 1326 -3757 1547 -3094
rect 2210 -3536 3315 -3315
rect 3978 -3536 4199 -3094
rect 1547 -3757 1768 -3315
rect 1989 -4420 2431 -3536
rect 1768 -3978 1989 -3536
rect 2431 -3757 2652 -3536
rect 3757 -3978 3978 -3315
rect 2873 -3757 3757 -3536
rect 3094 -3978 3757 -3757
rect 2431 -4420 3536 -3978
rect 1989 -4641 2210 -4420
rect 2431 -4641 2652 -4420
rect 2873 -4641 3094 -4420
rect 3315 -4641 3536 -4420
rect 663 -7514 884 -7293
rect 442 -7293 1105 -7072
rect 442 -7072 1326 -6851
rect 442 -6851 1768 -6630
rect 663 -6630 2210 -6409
rect 1768 -6409 2652 -6188
rect 2873 -6409 3757 -6188
rect 3315 -6630 5083 -6409
rect 3757 -6851 5083 -6630
rect 4199 -7072 5083 -6851
rect 4420 -7293 5083 -7072
rect 4641 -7514 4862 -7293
rect 2210 -6188 3315 -5746
rect 1768 -5746 2652 -5525
rect 2873 -5746 3757 -5525
rect 1326 -5525 2210 -5304
rect 3315 -5525 4199 -5304
rect 663 -5304 1989 -5083
rect 3536 -5304 4862 -5083
rect 442 -5083 1547 -4641
rect 3978 -5083 5083 -4641
rect 663 -4641 1326 -4420
rect 4199 -4641 4862 -4420
<< end >>
