magic
tech sky130A
magscale 1 2
timestamp 1735296899
<< metal1 >>
rect -756 12166 450 12266
rect 1884 12166 2930 12266
rect -4064 11998 -3246 12000
rect -756 11998 -656 12166
rect -4064 11900 -3116 11998
rect -7246 10692 -6572 10696
rect -4064 10692 -3964 11900
rect -3316 11898 -3116 11900
rect -1682 11898 -656 11998
rect 2830 11470 2930 12166
rect 2830 11370 3938 11470
rect 5372 11370 6150 11470
rect -7246 10596 -6444 10692
rect -7246 8462 -7146 10596
rect -6644 10592 -6444 10596
rect -5010 10592 -3964 10692
rect 6050 9680 6150 11370
rect 8562 9680 9368 9682
rect 6050 9580 7034 9680
rect 8468 9582 9368 9680
rect 8468 9580 8668 9582
rect -9722 8362 -9242 8462
rect -7808 8362 -7146 8462
rect -9722 5506 -9622 8362
rect 9268 7058 9368 9582
rect 9268 6958 9468 7058
rect 10902 7048 11102 7058
rect 10902 6958 11106 7048
rect 11006 6290 11106 6958
rect 11006 6190 12112 6290
rect -11456 5406 -11256 5506
rect -9822 5406 -9622 5506
rect -11456 3946 -11356 5406
rect -13052 3846 -11356 3946
rect -13052 2088 -12952 3846
rect 12012 3836 12112 6190
rect 10278 3828 10478 3836
rect 10276 3736 10478 3828
rect 11912 3736 12112 3836
rect -13052 1988 -12852 2088
rect -11418 2086 -11218 2088
rect -11418 1988 -10676 2086
rect -11384 1986 -10676 1988
rect -10776 -1488 -10676 1986
rect 10276 300 10376 3736
rect 10276 200 11554 300
rect 12988 280 13188 300
rect 12988 200 13190 280
rect -12510 -1588 -12310 -1488
rect -10876 -1588 -10676 -1488
rect -12510 -4910 -12410 -1588
rect 13090 -3236 13190 200
rect 10278 -3336 10478 -3236
rect 11912 -3336 13190 -3236
rect -11998 -4910 -11798 -4906
rect -12510 -5006 -11798 -4910
rect -10364 -4910 -10164 -4906
rect 10278 -4910 10378 -3336
rect -10364 -5006 -9884 -4910
rect -12510 -5010 -11958 -5006
rect -10330 -5010 -9884 -5006
rect 10278 -5010 10560 -4910
rect -9984 -8362 -9884 -5010
rect 10460 -6458 10560 -5010
rect 8388 -6558 8926 -6458
rect 10360 -6558 10560 -6458
rect -9984 -8462 -9784 -8362
rect -8350 -8462 -7846 -8362
rect -7946 -10596 -7846 -8462
rect 8388 -9580 8488 -6558
rect 6292 -9680 6492 -9580
rect 7926 -9680 8488 -9580
rect -7188 -10596 -6988 -10592
rect -7946 -10692 -6988 -10596
rect -5554 -10692 -4522 -10592
rect -7946 -10696 -7106 -10692
rect -4622 -11894 -4522 -10692
rect 3196 -11470 3396 -11370
rect 4830 -11376 5030 -11370
rect 6292 -11376 6392 -9680
rect 4830 -11470 6392 -11376
rect -4622 -11898 -3776 -11894
rect -4622 -11994 -3658 -11898
rect -3858 -11998 -3658 -11994
rect -2224 -11998 -1164 -11898
rect -1264 -12172 -1164 -11998
rect 3198 -12166 3298 -11470
rect 4918 -11476 6392 -11470
rect -292 -12172 -92 -12166
rect -1264 -12266 -92 -12172
rect 1342 -12266 3298 -12166
rect -1264 -12272 -212 -12266
<< metal2 >>
rect -199 14598 200 14600
rect -380 14595 380 14598
rect -561 14589 561 14595
rect -742 14581 742 14589
rect -923 14571 923 14581
rect -1104 14559 1104 14571
rect -1284 14544 1284 14559
rect -1465 14527 1465 14544
rect -1645 14508 1645 14527
rect -1825 14486 1825 14508
rect -2004 14462 2004 14486
rect -2184 14436 2184 14462
rect -2363 14408 2363 14436
rect -2541 14377 2541 14408
rect -2720 14344 2720 14377
rect -2898 14309 2898 14344
rect -3075 14272 3075 14309
rect -3252 14233 3252 14272
rect -3429 14198 3429 14233
rect -3429 14195 -161 14198
rect 161 14195 3429 14198
rect -3429 14191 -342 14195
rect -3605 14189 -342 14191
rect 342 14191 3429 14195
rect 342 14189 3605 14191
rect -3605 14181 -523 14189
rect 450 14181 3605 14189
rect -3605 14171 -704 14181
rect -3605 14159 -884 14171
rect -3605 14147 -1065 14159
rect -3781 14144 -1065 14147
rect -3781 14127 -1245 14144
rect -3781 14108 -1425 14127
rect -3781 14101 -1604 14108
rect -3956 14086 -1604 14101
rect -3956 14062 -1784 14086
rect -3956 14053 -1963 14062
rect -4130 14036 -1963 14053
rect -4130 14008 -2141 14036
rect -4130 14002 -2320 14008
rect -4304 13977 -2320 14002
rect -4304 13950 -2498 13977
rect -4477 13944 -2498 13950
rect -4477 13909 -2675 13944
rect -4477 13895 -2852 13909
rect -4649 13872 -2852 13895
rect -4649 13838 -3026 13872
rect -4821 13833 -3026 13838
rect -4821 13791 -3205 13833
rect -4821 13779 -3381 13791
rect -4992 13747 -3381 13779
rect -4992 13717 -3556 13747
rect -5162 13701 -3556 13717
rect -5162 13654 -3730 13701
rect -5332 13653 -3730 13654
rect -5332 13602 -3904 13653
rect -5332 13588 -4077 13602
rect -5500 13550 -4077 13588
rect -5500 13521 -4249 13550
rect -5668 13495 -4249 13521
rect -5668 13451 -4421 13495
rect -5835 13438 -4421 13451
rect -5835 13379 -4592 13438
rect -6001 13317 -4762 13379
rect -6001 13305 -4932 13317
rect -6167 13254 -4932 13305
rect -3116 13298 -3026 13833
rect 450 13566 540 14181
rect 704 14171 3605 14181
rect 884 14159 3605 14171
rect 1065 14147 3605 14159
rect 1065 14144 3781 14147
rect 1245 14127 3781 14144
rect 1425 14108 3781 14127
rect 1604 14101 3781 14108
rect 1604 14086 3956 14101
rect 1784 14062 3956 14086
rect 1963 14053 3956 14062
rect 1963 14036 4130 14053
rect 2141 14008 4130 14036
rect 2320 14002 4130 14008
rect 2320 13977 4304 14002
rect 2498 13950 4304 13977
rect 2498 13944 4477 13950
rect 2675 13909 4477 13944
rect 2852 13895 4477 13909
rect 2852 13872 4649 13895
rect 3029 13838 4649 13872
rect 3029 13833 4821 13838
rect 3205 13791 4821 13833
rect 3381 13779 4821 13791
rect 3381 13747 4992 13779
rect 3556 13717 4992 13747
rect 3556 13701 5162 13717
rect 3730 13654 5162 13701
rect 3730 13653 5332 13654
rect 3904 13602 5332 13653
rect -6167 13229 -5100 13254
rect -6331 13188 -5100 13229
rect -6331 13151 -5268 13188
rect -6494 13121 -5268 13151
rect -6494 13071 -5435 13121
rect -6656 13051 -5435 13071
rect -6656 12989 -5601 13051
rect -6817 12979 -5601 12989
rect -6817 12905 -5767 12979
rect -6817 12904 -5931 12905
rect -6978 12829 -5931 12904
rect -6978 12818 -6094 12829
rect -7137 12751 -6094 12818
rect 3938 12770 4028 13602
rect 4077 13588 5332 13602
rect 4077 13550 5500 13588
rect 4249 13521 5500 13550
rect 4249 13495 5668 13521
rect 4421 13451 5668 13495
rect 4421 13438 5835 13451
rect 4592 13379 5835 13438
rect 4762 13317 6001 13379
rect 4932 13305 6001 13317
rect 4932 13254 6167 13305
rect 5100 13229 6167 13254
rect 5100 13188 6331 13229
rect 5268 13151 6331 13188
rect 5268 13121 6494 13151
rect 5435 13071 6494 13121
rect 5435 13051 6656 13071
rect 5601 12989 6656 13051
rect 5601 12979 6817 12989
rect 5767 12905 6817 12979
rect 5931 12904 6817 12905
rect 5931 12829 6978 12904
rect 6094 12818 6978 12829
rect 6094 12751 7137 12818
rect -7137 12730 -6256 12751
rect -7295 12671 -6256 12730
rect 6256 12730 7137 12751
rect 6256 12671 7295 12730
rect -7295 12640 -6354 12671
rect -7452 12589 -6354 12640
rect 6417 12640 7295 12671
rect 6417 12589 7452 12640
rect -7452 12548 -6578 12589
rect -7607 12504 -6578 12548
rect -7607 12454 -6737 12504
rect -7762 12418 -6737 12454
rect -7762 12358 -6895 12418
rect -7915 12330 -6895 12358
rect -7915 12260 -7052 12330
rect -8068 12240 -7052 12260
rect -8068 12160 -7207 12240
rect -8219 12148 -7207 12160
rect -8219 12058 -7362 12148
rect -8368 12054 -7362 12058
rect -8368 11958 -7515 12054
rect -6444 11992 -6354 12589
rect 6578 12548 7452 12589
rect 6578 12504 7607 12548
rect 6737 12454 7607 12504
rect 6737 12418 7762 12454
rect 6895 12358 7762 12418
rect 6895 12330 7915 12358
rect 7034 12260 7915 12330
rect 7034 12240 8068 12260
rect -8368 11955 -7668 11958
rect -8517 11860 -7668 11955
rect -8517 11849 -7819 11860
rect -8664 11760 -7819 11849
rect -8664 11742 -7968 11760
rect -8809 11658 -7968 11742
rect -8809 11633 -8117 11658
rect -8954 11555 -8117 11633
rect -8954 11522 -8264 11555
rect -9097 11449 -8264 11522
rect -9097 11409 -8409 11449
rect -9238 11342 -8409 11409
rect -9238 11295 -8554 11342
rect -9378 11233 -8554 11295
rect -9378 11179 -8697 11233
rect -9517 11122 -8697 11179
rect -9517 11061 -8838 11122
rect -9654 11009 -8838 11061
rect -9654 10941 -8978 11009
rect 7034 10980 7124 12240
rect 7207 12160 8068 12240
rect 7207 12148 8219 12160
rect 7362 12058 8219 12148
rect 7362 12054 8368 12058
rect 7515 11958 8368 12054
rect 7668 11955 8368 11958
rect 7668 11860 8517 11955
rect 7819 11849 8517 11860
rect 7819 11760 8664 11849
rect 7968 11742 8664 11760
rect 7968 11658 8809 11742
rect 8117 11633 8809 11658
rect 8117 11555 8954 11633
rect 8264 11522 8954 11555
rect 8264 11449 9097 11522
rect 8409 11409 9097 11449
rect 8409 11342 9238 11409
rect 8554 11295 9238 11342
rect 8554 11233 9378 11295
rect 8697 11179 9378 11233
rect 8697 11122 9517 11179
rect 8838 11061 9517 11122
rect 8838 11009 9654 11061
rect -9790 10895 -8978 10941
rect 8978 10941 9654 11009
rect 8978 10895 9790 10941
rect -9790 10820 -9117 10895
rect -9924 10779 -9117 10820
rect 9117 10820 9790 10895
rect 9117 10779 9924 10820
rect -9924 10697 -9254 10779
rect -10057 10661 -9254 10697
rect -10057 10607 -9390 10661
rect -10057 10572 -9152 10607
rect -10188 10517 -9152 10572
rect -10188 10446 -9524 10517
rect -10318 10420 -9524 10446
rect -10318 10318 -9657 10420
rect -10446 10297 -9657 10318
rect -10446 10188 -9788 10297
rect -10572 10172 -9788 10188
rect -10572 10057 -9918 10172
rect -10697 10046 -9918 10057
rect -10697 9924 -10046 10046
rect -10820 9918 -10046 9924
rect -10820 9790 -10172 9918
rect -10941 9788 -10172 9790
rect -10941 9657 -10297 9788
rect -9242 9762 -9152 10517
rect -10941 9654 -10420 9657
rect -11061 9524 -10420 9654
rect -3116 9571 -3026 10498
rect -199 9998 200 10000
rect -371 9994 371 9998
rect 450 9994 540 10766
rect 9254 10697 9924 10779
rect 9254 10661 10057 10697
rect 9390 10572 10057 10661
rect 9390 10541 10188 10572
rect 9524 10446 10188 10541
rect 9524 10420 10318 10446
rect 9657 10318 10318 10420
rect 9657 10297 10446 10318
rect 9788 10188 10446 10297
rect 9788 10172 10572 10188
rect 9918 10057 10572 10172
rect 9918 10046 10697 10057
rect -542 9986 542 9994
rect -712 9976 712 9986
rect -883 9962 883 9976
rect -1054 9946 1054 9962
rect -1224 9926 1224 9946
rect -1394 9904 1394 9926
rect -1563 9879 1563 9904
rect -1733 9851 1733 9879
rect -1901 9819 1901 9851
rect -2069 9785 2069 9819
rect -2237 9748 2237 9785
rect -2404 9708 2404 9748
rect -2570 9666 2570 9708
rect -2736 9620 2736 9666
rect -2901 9598 2901 9620
rect -2901 9594 -142 9598
rect 142 9594 2901 9598
rect -2901 9586 -312 9594
rect 312 9586 2901 9594
rect -2901 9576 -483 9586
rect 483 9576 2901 9586
rect -2901 9571 -654 9576
rect -3116 9562 -654 9571
rect 654 9571 2901 9576
rect 654 9562 3065 9571
rect -3116 9546 -824 9562
rect 824 9546 3065 9562
rect -3116 9526 -994 9546
rect 994 9526 3065 9546
rect -11061 9517 -10541 9524
rect -3116 9520 -1163 9526
rect -11179 9390 -10541 9517
rect -3228 9504 -1163 9520
rect 1163 9520 3065 9526
rect 1163 9504 3228 9520
rect -3228 9479 -1333 9504
rect 1333 9479 3228 9504
rect -3228 9466 -1501 9479
rect -3390 9451 -1501 9466
rect 1501 9466 3228 9479
rect 1501 9451 3390 9466
rect -3390 9419 -1669 9451
rect 1669 9419 3390 9451
rect -3390 9408 -1837 9419
rect -11179 9378 -10661 9390
rect -11295 9254 -10661 9378
rect -3551 9385 -1837 9408
rect 1837 9408 3390 9419
rect 1837 9385 3551 9408
rect -3551 9349 -2004 9385
rect -3712 9348 -2004 9349
rect 2004 9349 3551 9385
rect 2004 9348 3712 9349
rect -3712 9308 -2170 9348
rect 2170 9308 3712 9348
rect -3712 9286 -2336 9308
rect -3871 9266 -2336 9286
rect 2336 9286 3712 9308
rect 2336 9266 3871 9286
rect -11295 9238 -10779 9254
rect -11409 9117 -10779 9238
rect -3871 9220 -2501 9266
rect 2501 9220 3871 9266
rect 3938 9220 4028 9970
rect 10046 9924 10697 10046
rect 10046 9918 10820 9924
rect 10172 9790 10820 9918
rect 10172 9788 10941 9790
rect 10297 9657 10941 9788
rect 10420 9654 10941 9657
rect 10420 9524 11061 9654
rect 10541 9517 11061 9524
rect 10541 9390 11179 9517
rect 10661 9378 11179 9390
rect 10661 9254 11295 9378
rect 10779 9238 11295 9254
rect -11409 9097 -10895 9117
rect -11522 8978 -10895 9097
rect -11522 8954 -11009 8978
rect -11633 8838 -11009 8954
rect -11633 8809 -11122 8838
rect -11742 8697 -11122 8809
rect -11742 8664 -11233 8697
rect -11849 8554 -11233 8664
rect -11849 8517 -11342 8554
rect -11955 8409 -11342 8517
rect -11955 8368 -11449 8409
rect -12058 8264 -11449 8368
rect -12058 8219 -11555 8264
rect -12160 8117 -11555 8219
rect -12160 8068 -11658 8117
rect -12260 7968 -11658 8068
rect -12260 7915 -11760 7968
rect -12358 7819 -11760 7915
rect -12358 7762 -11860 7819
rect -12454 7668 -11860 7762
rect -6444 7816 -6354 9192
rect -4029 9171 -2665 9220
rect 2665 9171 4029 9220
rect -4029 9152 -2828 9171
rect -4186 9120 -2828 9152
rect 2828 9152 4029 9171
rect 2828 9120 4186 9152
rect -4186 9081 -2990 9120
rect -4341 9066 -2990 9081
rect 2990 9081 4186 9120
rect 10779 9117 11409 9238
rect 10895 9097 11409 9117
rect 2990 9066 4341 9081
rect -4341 9008 -3151 9066
rect 3151 9008 4341 9066
rect -4496 8949 -3312 9008
rect 3312 8949 4496 9008
rect 10895 8978 11522 9097
rect -4496 8931 -3471 8949
rect -4649 8886 -3471 8931
rect 3471 8931 4496 8949
rect 11009 8954 11522 8978
rect 3471 8886 4649 8931
rect -4649 8852 -3629 8886
rect -4800 8820 -3629 8852
rect 3629 8852 4649 8886
rect 3629 8820 4800 8852
rect 11009 8838 11633 8954
rect -4800 8771 -3786 8820
rect -4951 8752 -3786 8771
rect 3786 8771 4800 8820
rect 11122 8809 11633 8838
rect 3786 8752 4951 8771
rect -4951 8687 -3941 8752
rect -5099 8681 -3941 8687
rect 3941 8687 4951 8752
rect 11122 8697 11742 8809
rect 3941 8681 5100 8687
rect -5099 8608 -4096 8681
rect 4096 8608 5100 8681
rect 11233 8664 11742 8697
rect 11233 8631 11849 8664
rect -5099 8600 -4249 8608
rect -5247 8531 -4249 8600
rect 4249 8600 5100 8608
rect 4249 8531 5247 8600
rect -5247 8510 -4400 8531
rect -5393 8452 -4400 8510
rect 4400 8510 5247 8531
rect 9468 8541 11849 8631
rect 4400 8452 5393 8510
rect -5393 8418 -4551 8452
rect -5537 8371 -4551 8418
rect 4551 8418 5393 8452
rect 4551 8371 5537 8418
rect -5537 8324 -4699 8371
rect -5680 8287 -4699 8324
rect 4700 8324 5537 8371
rect 9468 8358 9558 8541
rect 11342 8517 11849 8541
rect 11342 8409 11955 8517
rect 11449 8368 11955 8409
rect 4700 8287 5680 8324
rect -5680 8227 -4847 8287
rect -5821 8200 -4847 8227
rect 4847 8227 5680 8287
rect 11449 8264 12058 8368
rect 4847 8200 5821 8227
rect -5821 8128 -4993 8200
rect -5960 8110 -4993 8128
rect 4993 8128 5821 8200
rect 11555 8219 12058 8264
rect 4993 8110 5960 8128
rect -5960 8026 -5137 8110
rect -6097 8018 -5137 8026
rect 5137 8026 5960 8110
rect 5137 8018 6097 8026
rect -6097 7924 -5280 8018
rect 5280 7924 6097 8018
rect -6097 7922 -5421 7924
rect -6233 7827 -5421 7922
rect 5421 7922 6097 7924
rect 5421 7827 6233 7922
rect -6233 7816 -5560 7827
rect -6444 7728 -5560 7816
rect 5560 7816 6233 7827
rect 5560 7728 6367 7816
rect -6444 7707 -5697 7728
rect -12454 7607 -11958 7668
rect -12548 7515 -11958 7607
rect -6499 7626 -5697 7707
rect 5697 7707 6367 7728
rect 5697 7626 6499 7707
rect -6499 7596 -5833 7626
rect -6629 7522 -5833 7596
rect 5833 7596 6499 7626
rect 5833 7522 6629 7596
rect 7034 7529 7124 8180
rect 11555 8117 12160 8219
rect 11658 8068 12160 8117
rect 11658 7968 12260 8068
rect 11760 7915 12260 7968
rect 11760 7819 12358 7915
rect 11860 7762 12358 7819
rect 11860 7668 12454 7762
rect 11958 7607 12454 7668
rect -12548 7452 -12054 7515
rect -6629 7482 -5967 7522
rect -12640 7362 -12054 7452
rect -6757 7416 -5967 7482
rect 5967 7482 6629 7522
rect 5967 7416 6757 7482
rect -6757 7367 -6099 7416
rect -12640 7295 -12148 7362
rect -12730 7207 -12148 7295
rect -6883 7307 -6099 7367
rect 6099 7367 6757 7416
rect 6099 7307 6883 7367
rect -6883 7249 -6229 7307
rect -12730 7137 -12240 7207
rect -12818 7052 -12240 7137
rect -7007 7196 -6229 7249
rect 6229 7249 6883 7307
rect 7033 7249 7125 7529
rect 11958 7515 12548 7607
rect 12054 7452 12548 7515
rect 12054 7362 12640 7452
rect 6229 7196 7125 7249
rect 12148 7295 12640 7362
rect 12148 7207 12730 7295
rect -7007 7129 -6357 7196
rect -7129 7082 -6357 7129
rect 6357 7129 7125 7196
rect 12240 7137 12730 7207
rect 6357 7082 7129 7129
rect -12818 7006 -12330 7052
rect -7129 7007 -6483 7082
rect -12818 6978 -11166 7006
rect -12904 6916 -11166 6978
rect -7249 6967 -6483 7007
rect 6483 7007 7129 7082
rect 12240 7052 12818 7137
rect 6483 6967 7249 7007
rect -12904 6895 -12330 6916
rect -12904 6817 -12418 6895
rect -12989 6737 -12418 6817
rect -11256 6806 -11166 6916
rect -9242 6793 -9152 6962
rect -7249 6883 -6607 6967
rect -7367 6849 -6607 6883
rect 6607 6883 7249 6967
rect 12330 6978 12818 7052
rect 12330 6895 12904 6978
rect 6607 6849 7367 6883
rect -7367 6793 -6729 6849
rect -12989 6656 -12504 6737
rect -9242 6729 -6729 6793
rect 6729 6757 7367 6849
rect 12418 6817 12904 6895
rect 6729 6729 7482 6757
rect 12418 6737 12989 6817
rect -9242 6703 -6849 6729
rect -13071 6578 -12504 6656
rect -7482 6629 -6849 6703
rect -7596 6607 -6849 6629
rect 6849 6629 7482 6729
rect 12504 6656 12989 6737
rect 6849 6607 7596 6629
rect -13071 6494 -12589 6578
rect -7596 6499 -6967 6607
rect -13151 6417 -12589 6494
rect -7707 6483 -6967 6499
rect 6967 6499 7596 6607
rect 12504 6578 13071 6656
rect 6967 6483 7707 6499
rect -13151 6331 -12671 6417
rect -7707 6367 -7082 6483
rect -13229 6256 -12671 6331
rect -7816 6357 -7082 6367
rect 7082 6367 7707 6483
rect 12589 6494 13071 6578
rect 12589 6417 13151 6494
rect 7082 6357 7816 6367
rect -13229 6167 -12751 6256
rect -7816 6233 -7196 6357
rect -13305 6094 -12751 6167
rect -7922 6229 -7196 6233
rect 7196 6233 7816 6357
rect 12671 6331 13151 6417
rect 12671 6256 13229 6331
rect 7196 6229 7922 6233
rect -7922 6099 -7307 6229
rect 7307 6099 7922 6229
rect -7922 6097 -7416 6099
rect -13305 6001 -12829 6094
rect -13379 5931 -12829 6001
rect -8026 5967 -7416 6097
rect 7416 6097 7922 6099
rect 12751 6167 13229 6256
rect 7416 5967 8026 6097
rect 12751 6094 13305 6167
rect -8026 5960 -7522 5967
rect -13379 5835 -12905 5931
rect -13451 5767 -12905 5835
rect -8128 5833 -7522 5960
rect 7522 5960 8026 5967
rect 12829 6001 13305 6094
rect 7522 5833 8128 5960
rect 12829 5931 13379 6001
rect -8128 5821 -7626 5833
rect -13451 5668 -12979 5767
rect -8227 5697 -7626 5821
rect 7626 5821 8128 5833
rect 12905 5835 13379 5931
rect 7626 5697 8227 5821
rect 12905 5767 13451 5835
rect -8227 5680 -7728 5697
rect -13521 5601 -12979 5668
rect -13521 5500 -13051 5601
rect -8324 5560 -7728 5680
rect 7728 5680 8227 5697
rect 7728 5560 8324 5680
rect 12979 5668 13451 5767
rect 12979 5601 13521 5668
rect -8324 5537 -7827 5560
rect -13588 5435 -13051 5500
rect -13588 5332 -13121 5435
rect -8418 5421 -7827 5537
rect 7827 5537 8324 5560
rect 7827 5448 8418 5537
rect 9468 5448 9558 5558
rect 7827 5421 9558 5448
rect 13051 5500 13521 5601
rect 13051 5435 13588 5500
rect -8418 5393 -7924 5421
rect -13654 5268 -13121 5332
rect -8510 5280 -7924 5393
rect 7924 5358 9558 5421
rect 7924 5280 8510 5358
rect 13121 5336 13588 5435
rect -13654 5162 -13188 5268
rect -8510 5247 -8018 5280
rect -13717 5100 -13188 5162
rect -8600 5137 -8018 5247
rect 8018 5247 8510 5280
rect 11822 5332 13588 5336
rect 8018 5137 8600 5247
rect -13717 4992 -13254 5100
rect -8600 5099 -8110 5137
rect -13779 4932 -13254 4992
rect -8687 4993 -8110 5099
rect 8110 5099 8600 5137
rect 11822 5246 13654 5332
rect 11822 5136 11912 5246
rect 13188 5162 13654 5246
rect 13188 5100 13717 5162
rect 8110 4993 8687 5099
rect -8687 4951 -8200 4993
rect -13779 4821 -13317 4932
rect -13838 4762 -13317 4821
rect -8771 4847 -8200 4951
rect 8200 4951 8687 4993
rect 13254 4992 13717 5100
rect 8200 4847 8771 4951
rect 13254 4932 13779 4992
rect -8771 4800 -8287 4847
rect -13838 4649 -13379 4762
rect -8852 4699 -8287 4800
rect 8287 4800 8771 4847
rect 13317 4821 13779 4932
rect 8287 4699 8852 4800
rect 13317 4762 13838 4821
rect -8852 4649 -8371 4699
rect -13895 4592 -13379 4649
rect -13895 4477 -13438 4592
rect -8931 4551 -8371 4649
rect 8371 4649 8852 4699
rect 13379 4649 13838 4762
rect 8371 4551 8931 4649
rect 13379 4592 13895 4649
rect -8931 4496 -8452 4551
rect -13950 4421 -13438 4477
rect -13950 4304 -13495 4421
rect -9008 4400 -8452 4496
rect 8452 4496 8931 4551
rect 8452 4400 9008 4496
rect 13438 4477 13895 4592
rect 13438 4421 13950 4477
rect -9008 4341 -8531 4400
rect -14002 4249 -13495 4304
rect -9081 4249 -8531 4341
rect 8531 4341 9008 4400
rect 8531 4249 9081 4341
rect 13495 4304 13950 4421
rect 13495 4249 14002 4304
rect -14002 4130 -13550 4249
rect -9081 4186 -8608 4249
rect -14053 4077 -13550 4130
rect -9152 4096 -8608 4186
rect 8608 4186 9081 4249
rect 8608 4096 9152 4186
rect -14053 3956 -13602 4077
rect -9152 4029 -8681 4096
rect -14101 3904 -13602 3956
rect -14101 3781 -13653 3904
rect -11256 3896 -11166 4006
rect -9220 3941 -8681 4029
rect 8681 4029 9152 4096
rect 13550 4130 14002 4249
rect 13550 4077 14053 4130
rect 8681 3941 9220 4029
rect -9220 3896 -8752 3941
rect -11256 3806 -8752 3896
rect -14147 3730 -13653 3781
rect -9286 3786 -8752 3806
rect 8752 3871 9220 3941
rect 13602 3956 14053 4077
rect 13602 3904 14101 3956
rect 8752 3786 9286 3871
rect -14147 3605 -13701 3730
rect -9286 3712 -8820 3786
rect -14191 3579 -13701 3605
rect -9349 3629 -8820 3712
rect 8820 3712 9286 3786
rect 13653 3781 14101 3904
rect 13653 3730 14147 3781
rect 8820 3629 9349 3712
rect -11508 3579 -11418 3588
rect -14191 3489 -11418 3579
rect -9349 3551 -8886 3629
rect -14191 3429 -13747 3489
rect -14233 3381 -13747 3429
rect -11508 3388 -11418 3489
rect -9408 3471 -8886 3551
rect 8886 3551 9349 3629
rect 13701 3605 14147 3730
rect 13701 3556 14191 3605
rect 8886 3471 9408 3551
rect -9408 3390 -8949 3471
rect -14233 3252 -13791 3381
rect -14272 3205 -13791 3252
rect -9466 3312 -8949 3390
rect 8949 3390 9408 3471
rect 13747 3429 14191 3556
rect 8949 3312 9466 3390
rect 13747 3381 14233 3429
rect -9466 3228 -9008 3312
rect -14272 3075 -13833 3205
rect -14309 3029 -13833 3075
rect -9520 3151 -9008 3228
rect 9008 3228 9466 3312
rect 13791 3252 14233 3381
rect 9008 3151 9520 3228
rect 13791 3205 14272 3252
rect -9520 3065 -9066 3151
rect -14309 2898 -13872 3029
rect -9571 2990 -9066 3065
rect 9066 3065 9520 3151
rect 13833 3075 14272 3205
rect 9066 2990 9571 3065
rect 13833 3029 14309 3075
rect -9571 2901 -9120 2990
rect -14344 2852 -13872 2898
rect -14344 2720 -13909 2852
rect -9620 2828 -9120 2901
rect 9120 2901 9571 2990
rect 9120 2828 9620 2901
rect 13872 2898 14309 3029
rect 13872 2852 14344 2898
rect -9620 2736 -9171 2828
rect -14377 2675 -13909 2720
rect -14377 2541 -13944 2675
rect -9666 2665 -9171 2736
rect 9171 2736 9620 2828
rect 9171 2665 9666 2736
rect 13909 2720 14344 2852
rect 13909 2675 14377 2720
rect -9666 2570 -9220 2665
rect -14408 2498 -13944 2541
rect -9708 2501 -9220 2570
rect 9220 2570 9666 2665
rect 9220 2501 9708 2570
rect -14408 2363 -13977 2498
rect -9708 2404 -9266 2501
rect -14436 2320 -13977 2363
rect -9748 2336 -9266 2404
rect 9266 2404 9708 2501
rect 13944 2541 14377 2675
rect 13944 2498 14408 2541
rect 9266 2336 9748 2404
rect 13977 2363 14408 2498
rect -14436 2184 -14008 2320
rect -9748 2237 -9308 2336
rect -14462 2141 -14008 2184
rect -9785 2170 -9308 2237
rect 9308 2237 9748 2336
rect 9308 2226 9785 2237
rect 11822 2226 11912 2336
rect 13977 2320 14436 2363
rect 9308 2170 11912 2226
rect -14462 2004 -14036 2141
rect -9785 2069 -9348 2170
rect -14486 1963 -14036 2004
rect -9819 2004 -9348 2069
rect 9348 2136 11912 2170
rect 14008 2184 14436 2320
rect 14008 2141 14462 2184
rect 9348 2069 9785 2136
rect 9348 2004 9819 2069
rect -14486 1825 -14062 1963
rect -9819 1901 -9385 2004
rect -14508 1784 -14062 1825
rect -9851 1837 -9385 1901
rect 9385 1901 9819 2004
rect 14036 2004 14462 2141
rect 14036 1963 14486 2004
rect 9385 1837 9851 1901
rect -14508 1645 -14086 1784
rect -9851 1733 -9419 1837
rect -14527 1604 -14086 1645
rect -9879 1669 -9419 1733
rect 9419 1733 9851 1837
rect 14062 1825 14486 1963
rect 14062 1800 14508 1825
rect 9419 1669 9879 1733
rect -14527 1465 -14108 1604
rect -9879 1563 -9451 1669
rect -14544 1425 -14108 1465
rect -9904 1501 -9451 1563
rect 9451 1563 9879 1669
rect 11554 1710 14508 1800
rect 11554 1600 11644 1710
rect 14086 1645 14508 1710
rect 14086 1604 14527 1645
rect 9451 1501 9904 1563
rect -14544 1284 -14127 1425
rect -9904 1394 -9479 1501
rect -14559 1245 -14127 1284
rect -9926 1333 -9479 1394
rect 9479 1394 9904 1501
rect 14108 1465 14527 1604
rect 14108 1425 14544 1465
rect 9479 1333 9926 1394
rect -14559 1104 -14144 1245
rect -9926 1224 -9504 1333
rect -14571 1065 -14144 1104
rect -9946 1163 -9504 1224
rect 9504 1224 9926 1333
rect 14127 1284 14544 1425
rect 14127 1245 14559 1284
rect 9504 1163 9946 1224
rect -14571 923 -14159 1065
rect -9946 1054 -9526 1163
rect -14581 884 -14159 923
rect -9962 994 -9526 1054
rect 9526 1054 9946 1163
rect 14144 1104 14559 1245
rect 14144 1065 14571 1104
rect 9526 994 9962 1054
rect -14581 742 -14171 884
rect -9962 883 -9546 994
rect -14589 704 -14171 742
rect -9976 824 -9546 883
rect 9546 883 9962 994
rect 14159 923 14571 1065
rect 14159 884 14581 923
rect 9546 824 9976 883
rect -9976 712 -9562 824
rect -14589 561 -14181 704
rect -9986 654 -9562 712
rect 9562 712 9976 824
rect 14171 742 14581 884
rect 9562 654 9986 712
rect 14171 704 14589 742
rect -14595 523 -14181 561
rect -14595 380 -14189 523
rect -11508 487 -11418 588
rect -9986 542 -9576 654
rect -9994 487 -9576 542
rect -11508 483 -9576 487
rect 9576 542 9986 654
rect 14181 561 14589 704
rect 9576 483 9994 542
rect 14181 523 14595 561
rect -11508 397 -9586 483
rect -11508 388 -11418 397
rect -14598 342 -14189 380
rect -14598 200 -14195 342
rect -9998 312 -9586 397
rect 9586 371 9994 483
rect 14189 380 14595 523
rect 9586 312 9998 371
rect 14189 342 14598 380
rect -9998 200 -9594 312
rect -14600 161 -14195 200
rect -14600 12 -14198 161
rect -10000 142 -9594 200
rect 9594 200 9998 312
rect 14195 200 14598 342
rect 9594 142 10000 200
rect 14195 161 14600 200
rect -14600 -78 -12220 12
rect -14600 -161 -14198 -78
rect -14600 -199 -14195 -161
rect -12310 -188 -12220 -78
rect -10000 -142 -9598 142
rect 9598 -142 10000 142
rect -10000 -199 -9594 -142
rect -14598 -342 -14195 -199
rect -9998 -312 -9594 -199
rect 9594 -200 10000 -142
rect 14198 -161 14600 161
rect 14195 -200 14600 -161
rect 9594 -312 9998 -200
rect -14598 -380 -14189 -342
rect -9998 -371 -9586 -312
rect -14595 -523 -14189 -380
rect -9994 -483 -9586 -371
rect 9586 -371 9998 -312
rect 14195 -342 14598 -200
rect 9586 -483 9994 -371
rect -14595 -561 -14181 -523
rect -9994 -542 -9576 -483
rect -14589 -704 -14181 -561
rect -9986 -654 -9576 -542
rect 9576 -542 9994 -483
rect 14189 -380 14598 -342
rect 14189 -523 14595 -380
rect 9576 -654 9986 -542
rect -14589 -742 -14171 -704
rect -9986 -712 -9562 -654
rect -14581 -884 -14171 -742
rect -9976 -824 -9562 -712
rect 9562 -712 9986 -654
rect 14181 -561 14595 -523
rect 14181 -704 14589 -561
rect 9562 -824 9976 -712
rect -9976 -883 -9546 -824
rect -14581 -923 -14159 -884
rect -14571 -1065 -14159 -923
rect -9962 -994 -9546 -883
rect 9546 -883 9976 -824
rect 14171 -742 14589 -704
rect 9546 -994 9962 -883
rect 14171 -884 14581 -742
rect -9962 -1054 -9526 -994
rect -14571 -1104 -14144 -1065
rect -14559 -1245 -14144 -1104
rect -9946 -1163 -9526 -1054
rect 9526 -1054 9962 -994
rect 14159 -923 14581 -884
rect 9526 -1163 9946 -1054
rect 14159 -1065 14571 -923
rect -9946 -1224 -9504 -1163
rect -14559 -1284 -14127 -1245
rect -14544 -1425 -14127 -1284
rect -9926 -1333 -9504 -1224
rect 9504 -1224 9946 -1163
rect 14144 -1104 14571 -1065
rect 9504 -1310 9926 -1224
rect 11554 -1310 11644 -1200
rect 14144 -1245 14559 -1104
rect 9504 -1333 11644 -1310
rect -9926 -1394 -9479 -1333
rect -14544 -1465 -14108 -1425
rect -14527 -1604 -14108 -1465
rect -9904 -1501 -9479 -1394
rect 9479 -1400 11644 -1333
rect 14127 -1284 14559 -1245
rect 9479 -1501 9904 -1400
rect 14127 -1425 14544 -1284
rect -9904 -1563 -9451 -1501
rect -14527 -1645 -14086 -1604
rect -14508 -1784 -14086 -1645
rect -9879 -1669 -9451 -1563
rect 9451 -1563 9904 -1501
rect 14108 -1465 14544 -1425
rect 9451 -1669 9879 -1563
rect 14108 -1604 14527 -1465
rect -9879 -1733 -9419 -1669
rect -14508 -1825 -14062 -1784
rect -14486 -1963 -14062 -1825
rect -9851 -1837 -9419 -1733
rect 9419 -1733 9879 -1669
rect 14086 -1645 14527 -1604
rect 9419 -1837 9851 -1733
rect 14086 -1736 14508 -1645
rect -9851 -1901 -9385 -1837
rect -14486 -2004 -14036 -1963
rect -14462 -2141 -14036 -2004
rect -9819 -2004 -9385 -1901
rect 9385 -1901 9851 -1837
rect 11822 -1825 14508 -1736
rect 11822 -1826 14486 -1825
rect 9385 -2004 9819 -1901
rect 11822 -1936 11912 -1826
rect 14062 -1963 14486 -1826
rect -9819 -2069 -9348 -2004
rect -14462 -2184 -14008 -2141
rect -14436 -2320 -14008 -2184
rect -9785 -2170 -9348 -2069
rect 9348 -2069 9819 -2004
rect 14036 -2004 14486 -1963
rect 9348 -2170 9785 -2069
rect 14036 -2141 14462 -2004
rect -9785 -2237 -9308 -2170
rect -14436 -2363 -13977 -2320
rect -14408 -2498 -13977 -2363
rect -9748 -2336 -9308 -2237
rect 9308 -2237 9785 -2170
rect 14008 -2184 14462 -2141
rect 9308 -2336 9748 -2237
rect 14008 -2320 14436 -2184
rect -9748 -2404 -9266 -2336
rect -14408 -2541 -13944 -2498
rect -14377 -2675 -13944 -2541
rect -9708 -2501 -9266 -2404
rect 9266 -2404 9748 -2336
rect 13977 -2363 14436 -2320
rect 9266 -2501 9708 -2404
rect 13977 -2498 14408 -2363
rect -9708 -2570 -9220 -2501
rect -9666 -2665 -9220 -2570
rect 9220 -2570 9708 -2501
rect 13944 -2541 14408 -2498
rect 9220 -2665 9666 -2570
rect -14377 -2720 -13909 -2675
rect -14344 -2852 -13909 -2720
rect -9666 -2736 -9171 -2665
rect -9620 -2828 -9171 -2736
rect 9171 -2736 9666 -2665
rect 13944 -2675 14377 -2541
rect 13909 -2720 14377 -2675
rect 9171 -2828 9620 -2736
rect -14344 -2898 -13872 -2852
rect -14309 -3029 -13872 -2898
rect -9620 -2901 -9120 -2828
rect -14309 -3075 -13833 -3029
rect -14272 -3205 -13833 -3075
rect -12310 -3098 -12220 -2988
rect -9571 -2990 -9120 -2901
rect 9120 -2901 9620 -2828
rect 13909 -2852 14344 -2720
rect 13872 -2898 14344 -2852
rect 9120 -2990 9571 -2901
rect -9571 -3065 -9066 -2990
rect -9520 -3098 -9066 -3065
rect -12310 -3151 -9066 -3098
rect 9066 -3065 9571 -2990
rect 13872 -3029 14309 -2898
rect 9066 -3151 9520 -3065
rect -12310 -3188 -9008 -3151
rect -14272 -3252 -13791 -3205
rect -9520 -3228 -9008 -3188
rect -14233 -3381 -13791 -3252
rect -9466 -3312 -9008 -3228
rect 9008 -3228 9520 -3151
rect 13833 -3075 14309 -3029
rect 13833 -3205 14272 -3075
rect 9008 -3312 9466 -3228
rect -14233 -3406 -13747 -3381
rect -9466 -3390 -8949 -3312
rect -14233 -3429 -10364 -3406
rect -14191 -3496 -10364 -3429
rect -14191 -3556 -13747 -3496
rect -14191 -3605 -13701 -3556
rect -14147 -3730 -13701 -3605
rect -10454 -3606 -10364 -3496
rect -9408 -3471 -8949 -3390
rect 8949 -3390 9466 -3312
rect 13791 -3252 14272 -3205
rect 13791 -3381 14233 -3252
rect 8949 -3471 9408 -3390
rect -9408 -3551 -8886 -3471
rect -9349 -3629 -8886 -3551
rect 8886 -3551 9408 -3471
rect 13747 -3429 14233 -3381
rect 8886 -3629 9349 -3551
rect 13747 -3556 14191 -3429
rect -9349 -3712 -8820 -3629
rect -14147 -3781 -13653 -3730
rect -14101 -3904 -13653 -3781
rect -9286 -3786 -8820 -3712
rect 8820 -3712 9349 -3629
rect 13701 -3605 14191 -3556
rect 8820 -3786 9286 -3712
rect 13701 -3730 14147 -3605
rect -9286 -3871 -8752 -3786
rect -14101 -3956 -13602 -3904
rect -14053 -4077 -13602 -3956
rect -9220 -3941 -8752 -3871
rect 8752 -3871 9286 -3786
rect 13653 -3781 14147 -3730
rect 8752 -3941 9220 -3871
rect 13653 -3904 14101 -3781
rect -9220 -4029 -8681 -3941
rect -14053 -4130 -13550 -4077
rect -14002 -4249 -13550 -4130
rect -9152 -4096 -8681 -4029
rect 8681 -4029 9220 -3941
rect 13602 -3956 14101 -3904
rect 8681 -4096 9152 -4029
rect 13602 -4077 14053 -3956
rect -9152 -4186 -8608 -4096
rect -9081 -4249 -8608 -4186
rect 8608 -4186 9152 -4096
rect 13550 -4130 14053 -4077
rect 8608 -4249 9081 -4186
rect 13550 -4249 14002 -4130
rect -14002 -4304 -13495 -4249
rect -13950 -4421 -13495 -4304
rect -9081 -4341 -8531 -4249
rect -9008 -4400 -8531 -4341
rect 8531 -4341 9081 -4249
rect 13495 -4304 14002 -4249
rect 8531 -4400 9008 -4341
rect -13950 -4477 -13438 -4421
rect -13895 -4592 -13438 -4477
rect -9008 -4496 -8452 -4400
rect -8931 -4551 -8452 -4496
rect 8452 -4496 9008 -4400
rect 13495 -4421 13950 -4304
rect 13438 -4477 13950 -4421
rect 8452 -4551 8931 -4496
rect -13895 -4649 -13379 -4592
rect -8931 -4649 -8371 -4551
rect -13838 -4762 -13379 -4649
rect -8852 -4700 -8371 -4649
rect 8371 -4649 8931 -4551
rect 13438 -4592 13895 -4477
rect 13379 -4649 13895 -4592
rect 8371 -4700 8852 -4649
rect -13838 -4821 -13317 -4762
rect -8852 -4800 -8287 -4700
rect -13779 -4932 -13317 -4821
rect -8771 -4847 -8287 -4800
rect 8287 -4800 8852 -4700
rect 8287 -4846 8771 -4800
rect 11822 -4846 11912 -4736
rect 13379 -4762 13838 -4649
rect 8287 -4847 11912 -4846
rect -13779 -4992 -13254 -4932
rect -8771 -4951 -8200 -4847
rect -13717 -5100 -13254 -4992
rect -8687 -4993 -8200 -4951
rect 8200 -4936 11912 -4847
rect 13317 -4821 13838 -4762
rect 13317 -4932 13779 -4821
rect 8200 -4951 8771 -4936
rect 8200 -4993 8687 -4951
rect -8687 -5100 -8110 -4993
rect -13717 -5162 -13188 -5100
rect -13654 -5268 -13188 -5162
rect -8600 -5137 -8110 -5100
rect 8110 -5100 8687 -4993
rect 13254 -4992 13779 -4932
rect 13254 -5015 13717 -4992
rect 8110 -5137 8600 -5100
rect -8600 -5247 -8018 -5137
rect -13654 -5332 -13121 -5268
rect -13588 -5435 -13121 -5332
rect -8510 -5280 -8018 -5247
rect 8018 -5247 8600 -5137
rect 10270 -5105 13717 -5015
rect 10270 -5158 10360 -5105
rect 13188 -5162 13717 -5105
rect 8018 -5280 8510 -5247
rect 13188 -5268 13654 -5162
rect -8510 -5393 -7924 -5280
rect -8418 -5421 -7924 -5393
rect 7924 -5393 8510 -5280
rect 13121 -5332 13654 -5268
rect 7924 -5421 8418 -5393
rect -13588 -5500 -13051 -5435
rect -13521 -5601 -13051 -5500
rect -8418 -5537 -7827 -5421
rect -8324 -5560 -7827 -5537
rect 7827 -5537 8418 -5421
rect 13121 -5435 13588 -5332
rect 13051 -5500 13588 -5435
rect 7827 -5560 8324 -5537
rect -13521 -5668 -12979 -5601
rect -13451 -5767 -12979 -5668
rect -8324 -5680 -7728 -5560
rect -8227 -5697 -7728 -5680
rect 7728 -5680 8324 -5560
rect 13051 -5601 13521 -5500
rect 12979 -5668 13521 -5601
rect 7728 -5697 8227 -5680
rect -13451 -5835 -12905 -5767
rect -8227 -5821 -7626 -5697
rect -13379 -5931 -12905 -5835
rect -8128 -5833 -7626 -5821
rect 7626 -5821 8227 -5697
rect 12979 -5767 13451 -5668
rect 7626 -5833 8128 -5821
rect -13379 -6001 -12829 -5931
rect -8128 -5960 -7522 -5833
rect -13305 -6094 -12829 -6001
rect -8026 -5967 -7522 -5960
rect 7522 -5960 8128 -5833
rect 12905 -5835 13451 -5767
rect 12905 -5931 13379 -5835
rect 7522 -5967 8026 -5960
rect -13305 -6167 -12751 -6094
rect -8026 -6097 -7416 -5967
rect -13229 -6256 -12751 -6167
rect -7922 -6099 -7416 -6097
rect 7416 -6097 8026 -5967
rect 12829 -6001 13379 -5931
rect 12829 -6094 13305 -6001
rect 7416 -6099 7922 -6097
rect -7922 -6229 -7307 -6099
rect 7307 -6229 7922 -6099
rect -7922 -6233 -7196 -6229
rect -13229 -6331 -12671 -6256
rect -13151 -6417 -12671 -6331
rect -7841 -6357 -7196 -6233
rect 7196 -6233 7922 -6229
rect 12751 -6167 13305 -6094
rect 7196 -6357 7816 -6233
rect 12751 -6256 13229 -6167
rect -7841 -6367 -7082 -6357
rect -13151 -6494 -12589 -6417
rect -13071 -6578 -12589 -6494
rect -10454 -6516 -10364 -6406
rect -7841 -6516 -7751 -6367
rect -7707 -6483 -7082 -6367
rect 7082 -6367 7816 -6357
rect 12671 -6331 13229 -6256
rect 7082 -6483 7707 -6367
rect 12671 -6417 13151 -6331
rect -7707 -6499 -6967 -6483
rect -13071 -6656 -12504 -6578
rect -10454 -6606 -7751 -6516
rect -7596 -6607 -6967 -6499
rect 6967 -6499 7707 -6483
rect 12589 -6494 13151 -6417
rect 6967 -6607 7596 -6499
rect 12589 -6578 13071 -6494
rect -7596 -6629 -6849 -6607
rect -12989 -6737 -12504 -6656
rect -7482 -6673 -6849 -6629
rect -8440 -6729 -6849 -6673
rect 6849 -6629 7596 -6607
rect 6849 -6729 7482 -6629
rect -12989 -6817 -12418 -6737
rect -12904 -6895 -12418 -6817
rect -8440 -6763 -6729 -6729
rect -12904 -6978 -12330 -6895
rect -8440 -6962 -8350 -6763
rect -7367 -6849 -6729 -6763
rect 6729 -6757 7482 -6729
rect 12504 -6656 13071 -6578
rect 12504 -6737 12989 -6656
rect 6729 -6849 7367 -6757
rect -7367 -6883 -6607 -6849
rect -12818 -7052 -12330 -6978
rect -7249 -6967 -6607 -6883
rect 6607 -6883 7367 -6849
rect 12418 -6817 12989 -6737
rect 6607 -6967 7249 -6883
rect 12418 -6895 12904 -6817
rect -7249 -7007 -6483 -6967
rect -12818 -7137 -12240 -7052
rect -7129 -7082 -6483 -7007
rect 6483 -7007 7249 -6967
rect 12330 -6978 12904 -6895
rect 6483 -7082 7129 -7007
rect 12330 -7052 12818 -6978
rect -7129 -7129 -6357 -7082
rect -12730 -7207 -12240 -7137
rect -7007 -7196 -6357 -7129
rect 6357 -7129 7129 -7082
rect 6357 -7196 7007 -7129
rect -12730 -7295 -12148 -7207
rect -7007 -7249 -6229 -7196
rect -12640 -7362 -12148 -7295
rect -6883 -7307 -6229 -7249
rect 6229 -7249 7007 -7196
rect 12240 -7137 12818 -7052
rect 12240 -7207 12730 -7137
rect 6229 -7307 6883 -7249
rect -12640 -7452 -12054 -7362
rect -6883 -7367 -6099 -7307
rect -12548 -7515 -12054 -7452
rect -6757 -7416 -6099 -7367
rect 6099 -7367 6883 -7307
rect 12148 -7295 12730 -7207
rect 12148 -7362 12640 -7295
rect 6099 -7416 6757 -7367
rect -6757 -7482 -5967 -7416
rect -12548 -7607 -11958 -7515
rect -6629 -7522 -5967 -7482
rect 5967 -7482 6757 -7416
rect 12054 -7452 12640 -7362
rect 5967 -7522 6629 -7482
rect 12054 -7515 12548 -7452
rect -6629 -7596 -5833 -7522
rect -12454 -7668 -11958 -7607
rect -6499 -7626 -5833 -7596
rect 5833 -7596 6629 -7522
rect 5833 -7626 6499 -7596
rect -12454 -7762 -11860 -7668
rect -6499 -7707 -5697 -7626
rect -12358 -7819 -11860 -7762
rect -6367 -7728 -5697 -7707
rect 5697 -7707 6499 -7626
rect 11958 -7607 12548 -7515
rect 11958 -7668 12454 -7607
rect 5697 -7728 6367 -7707
rect -6367 -7816 -5560 -7728
rect -12358 -7915 -11760 -7819
rect -12260 -7968 -11760 -7915
rect -6233 -7827 -5560 -7816
rect 5560 -7816 6367 -7728
rect 11860 -7762 12454 -7668
rect 5560 -7827 6233 -7816
rect 11860 -7819 12358 -7762
rect -6233 -7922 -5421 -7827
rect -6097 -7924 -5421 -7922
rect 5421 -7922 6233 -7827
rect 11760 -7915 12358 -7819
rect 5421 -7924 6097 -7922
rect -12260 -8068 -11658 -7968
rect -6097 -8018 -5280 -7924
rect 5280 -8018 6097 -7924
rect -6097 -8026 -5137 -8018
rect -12160 -8117 -11658 -8068
rect -5960 -8110 -5137 -8026
rect 5137 -8026 6097 -8018
rect 5137 -8068 5960 -8026
rect 10270 -8068 10360 -7958
rect 11760 -7968 12260 -7915
rect 5137 -8110 10360 -8068
rect -12160 -8219 -11555 -8117
rect -5960 -8128 -4993 -8110
rect -12058 -8264 -11555 -8219
rect -5821 -8200 -4993 -8128
rect 4993 -8158 10360 -8110
rect 11658 -8068 12260 -7968
rect 11658 -8117 12160 -8068
rect 4993 -8200 5821 -8158
rect 7836 -8180 7926 -8158
rect -5821 -8227 -4847 -8200
rect -12058 -8368 -11449 -8264
rect -5680 -8287 -4847 -8227
rect 4847 -8227 5821 -8200
rect 11555 -8219 12160 -8117
rect 4847 -8287 5680 -8227
rect 11555 -8264 12058 -8219
rect -5680 -8324 -4700 -8287
rect -11955 -8409 -11449 -8368
rect -5644 -8371 -4700 -8324
rect 4700 -8324 5680 -8287
rect 4700 -8371 5537 -8324
rect -11955 -8517 -11342 -8409
rect -11849 -8554 -11342 -8517
rect -5644 -8418 -4551 -8371
rect -11849 -8664 -11233 -8554
rect -11742 -8697 -11233 -8664
rect -11742 -8809 -11122 -8697
rect -11633 -8838 -11122 -8809
rect -11633 -8954 -11009 -8838
rect -11522 -8978 -11009 -8954
rect -11522 -9097 -10895 -8978
rect -11409 -9117 -10895 -9097
rect -11409 -9238 -10779 -9117
rect -5644 -9192 -5554 -8418
rect -5393 -8452 -4551 -8418
rect 4551 -8418 5537 -8371
rect 11449 -8368 12058 -8264
rect 11449 -8409 11955 -8368
rect 4551 -8452 5393 -8418
rect -5393 -8510 -4400 -8452
rect -5247 -8531 -4400 -8510
rect 4400 -8510 5393 -8452
rect 4400 -8531 5247 -8510
rect -5247 -8600 -4249 -8531
rect -5100 -8608 -4249 -8600
rect 4249 -8600 5247 -8531
rect 11342 -8517 11955 -8409
rect 11342 -8554 11849 -8517
rect 4249 -8608 5100 -8600
rect -5100 -8681 -4096 -8608
rect 4096 -8681 5100 -8608
rect -5100 -8687 -3941 -8681
rect -4951 -8752 -3941 -8687
rect 3941 -8687 5100 -8681
rect 11233 -8664 11849 -8554
rect 3941 -8752 4951 -8687
rect 11233 -8697 11742 -8664
rect -4951 -8771 -3786 -8752
rect -4800 -8820 -3786 -8771
rect 3786 -8771 4951 -8752
rect 3786 -8820 4830 -8771
rect -4800 -8852 -3629 -8820
rect -4649 -8886 -3629 -8852
rect 3629 -8852 4830 -8820
rect 11122 -8809 11742 -8697
rect 11122 -8838 11633 -8809
rect 3629 -8886 4649 -8852
rect -4649 -8931 -3471 -8886
rect -4496 -8949 -3471 -8931
rect 3471 -8931 4649 -8886
rect 3471 -8949 4496 -8931
rect -4496 -9008 -3312 -8949
rect 3312 -9008 4496 -8949
rect -4341 -9066 -3151 -9008
rect 3151 -9066 4341 -9008
rect -4341 -9081 -2990 -9066
rect -4186 -9120 -2990 -9081
rect 2990 -9081 4341 -9066
rect 2990 -9120 4186 -9081
rect -4186 -9152 -2828 -9120
rect -4029 -9171 -2828 -9152
rect 2828 -9152 4186 -9120
rect 2828 -9171 4029 -9152
rect -4029 -9220 -2665 -9171
rect 2665 -9220 4029 -9171
rect -11295 -9254 -10779 -9238
rect -11295 -9378 -10661 -9254
rect -3871 -9266 -2501 -9220
rect 2501 -9266 3871 -9220
rect -3871 -9286 -2336 -9266
rect -3712 -9308 -2336 -9286
rect 2336 -9286 3871 -9266
rect 2336 -9308 3712 -9286
rect -3712 -9348 -2170 -9308
rect 2170 -9348 3712 -9308
rect -3712 -9349 -2004 -9348
rect -11179 -9390 -10661 -9378
rect -3551 -9385 -2004 -9349
rect 2004 -9349 3712 -9348
rect 2004 -9385 3551 -9349
rect -11179 -9517 -10541 -9390
rect -3551 -9408 -1837 -9385
rect -3390 -9419 -1837 -9408
rect 1837 -9408 3551 -9385
rect 1837 -9419 3390 -9408
rect -3390 -9451 -1669 -9419
rect 1669 -9451 3390 -9419
rect -3390 -9466 -1501 -9451
rect -11061 -9524 -10541 -9517
rect -3228 -9479 -1501 -9466
rect 1501 -9466 3390 -9451
rect 1501 -9479 3228 -9466
rect -3228 -9504 -1333 -9479
rect 1333 -9504 3228 -9479
rect -3228 -9520 -1163 -9504
rect -11061 -9654 -10420 -9524
rect -3065 -9526 -1163 -9520
rect 1163 -9520 3228 -9504
rect 1163 -9526 3065 -9520
rect -3065 -9546 -994 -9526
rect 994 -9546 3065 -9526
rect -3065 -9562 -824 -9546
rect 824 -9562 3065 -9546
rect -3065 -9571 -654 -9562
rect -2901 -9576 -654 -9571
rect 654 -9571 3065 -9562
rect 654 -9576 2901 -9571
rect -2901 -9586 -483 -9576
rect 483 -9586 2901 -9576
rect -2901 -9594 -312 -9586
rect 312 -9594 2901 -9586
rect -2901 -9598 -142 -9594
rect 142 -9598 2901 -9594
rect -2901 -9620 2901 -9598
rect -10941 -9657 -10420 -9654
rect -10941 -9788 -10297 -9657
rect -2736 -9666 2736 -9620
rect -2570 -9708 2570 -9666
rect -2404 -9748 2404 -9708
rect -10941 -9790 -10172 -9788
rect -10820 -9918 -10172 -9790
rect -10820 -9924 -10046 -9918
rect -10697 -10046 -10046 -9924
rect -10697 -10057 -9918 -10046
rect -10572 -10172 -9918 -10057
rect -10572 -10188 -9788 -10172
rect -10446 -10297 -9788 -10188
rect -10446 -10318 -9657 -10297
rect -10318 -10420 -9657 -10318
rect -10318 -10446 -9524 -10420
rect -10188 -10541 -9524 -10446
rect -10188 -10572 -9390 -10541
rect -10057 -10661 -9390 -10572
rect -10057 -10697 -9254 -10661
rect -9924 -10779 -9254 -10697
rect -9924 -10820 -9117 -10779
rect -9790 -10895 -9117 -10820
rect -9790 -10941 -8978 -10895
rect -9654 -11009 -8978 -10941
rect -9654 -11061 -8838 -11009
rect -9517 -11122 -8838 -11061
rect -9517 -11179 -8697 -11122
rect -9378 -11233 -8697 -11179
rect -9378 -11295 -8554 -11233
rect -9238 -11342 -8554 -11295
rect -8440 -11342 -8350 -9762
rect -2314 -9785 2237 -9748
rect -2314 -10498 -2224 -9785
rect -2069 -9819 2069 -9785
rect -1901 -9851 1901 -9819
rect -1733 -9879 1733 -9851
rect -1563 -9904 1563 -9879
rect -1394 -9926 1394 -9904
rect -1224 -9946 1224 -9926
rect -1054 -9962 1054 -9946
rect -883 -9976 883 -9962
rect -712 -9986 712 -9976
rect -542 -9994 542 -9986
rect -371 -9998 371 -9994
rect -200 -10000 199 -9998
rect 1252 -10766 1342 -9926
rect 4740 -9970 4830 -8852
rect 11009 -8954 11633 -8838
rect 11009 -8978 11522 -8954
rect 10895 -9097 11522 -8978
rect 10895 -9117 11409 -9097
rect 10779 -9238 11409 -9117
rect 10779 -9254 11295 -9238
rect 10661 -9378 11295 -9254
rect 10661 -9390 11179 -9378
rect 10541 -9517 11179 -9390
rect 10541 -9524 11061 -9517
rect 10420 -9654 11061 -9524
rect 10420 -9657 10941 -9654
rect 10297 -9788 10941 -9657
rect 10172 -9790 10941 -9788
rect 10172 -9918 10820 -9790
rect 10046 -9924 10820 -9918
rect 10046 -10046 10697 -9924
rect 9918 -10057 10697 -10046
rect 9918 -10172 10572 -10057
rect 9788 -10188 10572 -10172
rect 9788 -10297 10446 -10188
rect 9657 -10318 10446 -10297
rect 9657 -10420 10318 -10318
rect 9524 -10446 10318 -10420
rect 9524 -10541 10188 -10446
rect 9390 -10572 10188 -10541
rect 9390 -10661 10057 -10572
rect 9254 -10697 10057 -10661
rect 9254 -10779 9924 -10697
rect 9117 -10820 9924 -10779
rect 9117 -10895 9790 -10820
rect 8978 -10941 9790 -10895
rect 7836 -11090 7926 -10980
rect 8978 -11009 9654 -10941
rect 8838 -11061 9654 -11009
rect 8838 -11090 9517 -11061
rect 7836 -11179 9517 -11090
rect 7836 -11180 9378 -11179
rect 8697 -11233 9378 -11180
rect 8554 -11295 9378 -11233
rect 8554 -11342 9238 -11295
rect -9238 -11409 -8350 -11342
rect -9097 -11449 -8350 -11409
rect 8409 -11409 9238 -11342
rect 8409 -11449 9097 -11409
rect -9097 -11522 -8264 -11449
rect -8954 -11555 -8264 -11522
rect 8264 -11522 9097 -11449
rect 8264 -11555 8954 -11522
rect -8954 -11633 -8117 -11555
rect -8809 -11658 -8117 -11633
rect 8117 -11633 8954 -11555
rect 8117 -11658 8809 -11633
rect -8809 -11742 -7968 -11658
rect -8664 -11760 -7968 -11742
rect 7968 -11742 8809 -11658
rect 7968 -11760 8664 -11742
rect -8664 -11849 -7819 -11760
rect -8517 -11860 -7819 -11849
rect 7819 -11849 8664 -11760
rect 7819 -11860 8517 -11849
rect -8517 -11955 -7668 -11860
rect -8368 -11958 -7668 -11955
rect 7668 -11955 8517 -11860
rect 7668 -11958 8368 -11955
rect -8368 -12054 -7515 -11958
rect -8368 -12058 -7362 -12054
rect -8219 -12148 -7362 -12058
rect -8219 -12160 -7207 -12148
rect -8068 -12240 -7207 -12160
rect -8068 -12260 -7052 -12240
rect -7915 -12330 -7052 -12260
rect -7915 -12358 -6895 -12330
rect -7762 -12418 -6895 -12358
rect -7762 -12454 -6737 -12418
rect -7607 -12504 -6737 -12454
rect -7607 -12548 -6578 -12504
rect -7452 -12589 -6578 -12548
rect -7452 -12640 -6417 -12589
rect -7295 -12671 -6417 -12640
rect -7295 -12730 -6256 -12671
rect -7137 -12751 -6256 -12730
rect -7137 -12818 -6094 -12751
rect -6978 -12829 -6094 -12818
rect -6978 -12904 -5931 -12829
rect -6817 -12905 -5931 -12904
rect -6817 -12979 -5767 -12905
rect -5644 -12979 -5554 -11992
rect 7515 -12054 8368 -11958
rect 7362 -12058 8368 -12054
rect 7362 -12148 8219 -12058
rect 7207 -12160 8219 -12148
rect 7207 -12240 8068 -12160
rect 7052 -12260 8068 -12240
rect 7052 -12330 7915 -12260
rect 6895 -12358 7915 -12330
rect 6895 -12418 7762 -12358
rect 6737 -12454 7762 -12418
rect 6737 -12504 7607 -12454
rect 6578 -12548 7607 -12504
rect 6578 -12589 7452 -12548
rect 6417 -12640 7452 -12589
rect 6417 -12671 7295 -12640
rect 6256 -12730 7295 -12671
rect 6256 -12751 7137 -12730
rect -6817 -12989 -5554 -12979
rect -6656 -13051 -5554 -12989
rect -6656 -13071 -5435 -13051
rect -6494 -13121 -5435 -13071
rect -6494 -13151 -5268 -13121
rect -6331 -13188 -5268 -13151
rect -6331 -13229 -5100 -13188
rect -6167 -13254 -5100 -13229
rect -6167 -13305 -4932 -13254
rect -6001 -13317 -4932 -13305
rect -6001 -13379 -4762 -13317
rect -5835 -13438 -4592 -13379
rect -5835 -13451 -4421 -13438
rect -5668 -13495 -4421 -13451
rect -5668 -13521 -4249 -13495
rect -2314 -13515 -2224 -13298
rect 4740 -13317 4830 -12770
rect 6094 -12818 7137 -12751
rect 6094 -12829 6978 -12818
rect 5931 -12904 6978 -12829
rect 5931 -12905 6817 -12904
rect 5767 -12979 6817 -12905
rect 5601 -12989 6817 -12979
rect 5601 -13051 6656 -12989
rect 5435 -13071 6656 -13051
rect 5435 -13121 6494 -13071
rect 5268 -13151 6494 -13121
rect 5268 -13188 6331 -13151
rect 5100 -13229 6331 -13188
rect 5100 -13254 6167 -13229
rect 4932 -13305 6167 -13254
rect 4932 -13317 6001 -13305
rect 4740 -13379 6001 -13317
rect 4592 -13438 5835 -13379
rect 4421 -13451 5835 -13438
rect 4421 -13495 5668 -13451
rect -5500 -13550 -4249 -13521
rect -5500 -13588 -4077 -13550
rect -5332 -13602 -4077 -13588
rect -5332 -13653 -3904 -13602
rect -2377 -13605 -2224 -13515
rect 4249 -13521 5668 -13495
rect 4249 -13550 5500 -13521
rect -5332 -13654 -3730 -13653
rect -5162 -13701 -3730 -13654
rect -5162 -13717 -3556 -13701
rect -4992 -13747 -3556 -13717
rect -4992 -13779 -3381 -13747
rect -4821 -13791 -3381 -13779
rect -4821 -13833 -3205 -13791
rect -4821 -13838 -3029 -13833
rect -4649 -13872 -3029 -13838
rect -4649 -13895 -2852 -13872
rect -4477 -13909 -2852 -13895
rect -4477 -13944 -2675 -13909
rect -4477 -13950 -2498 -13944
rect -4304 -13977 -2498 -13950
rect -2377 -13977 -2287 -13605
rect -4304 -14002 -2287 -13977
rect -4130 -14008 -2287 -14002
rect -4130 -14036 -2141 -14008
rect -4130 -14053 -1963 -14036
rect -3956 -14062 -1963 -14053
rect -3956 -14086 -1784 -14062
rect -3956 -14101 -1604 -14086
rect -3781 -14108 -1604 -14101
rect -3781 -14127 -1425 -14108
rect 1252 -14127 1342 -13566
rect 4077 -13588 5500 -13550
rect 4077 -13602 5332 -13588
rect 3904 -13653 5332 -13602
rect 3730 -13654 5332 -13653
rect 3730 -13701 5162 -13654
rect 3556 -13717 5162 -13701
rect 3556 -13747 4992 -13717
rect 3381 -13779 4992 -13747
rect 3381 -13791 4821 -13779
rect 3205 -13833 4821 -13791
rect 3029 -13838 4821 -13833
rect 3029 -13872 4649 -13838
rect 2852 -13895 4649 -13872
rect 2852 -13909 4477 -13895
rect 2675 -13944 4477 -13909
rect 2498 -13950 4477 -13944
rect 2498 -13977 4304 -13950
rect 2320 -14002 4304 -13977
rect 2320 -14008 4130 -14002
rect 2141 -14036 4130 -14008
rect 1963 -14053 4130 -14036
rect 1963 -14062 3956 -14053
rect 1784 -14086 3956 -14062
rect 1604 -14101 3956 -14086
rect 1604 -14108 3781 -14101
rect 1425 -14127 3781 -14108
rect -3781 -14144 -1245 -14127
rect 1245 -14144 3781 -14127
rect -3781 -14147 -1065 -14144
rect -3605 -14159 -1065 -14147
rect 1065 -14147 3781 -14144
rect 1065 -14159 3605 -14147
rect -3605 -14171 -884 -14159
rect 884 -14171 3605 -14159
rect -3605 -14181 -704 -14171
rect 704 -14181 3605 -14171
rect -3605 -14189 -523 -14181
rect 523 -14189 3605 -14181
rect -3605 -14191 -342 -14189
rect -3429 -14195 -342 -14191
rect 342 -14191 3605 -14189
rect 342 -14195 3429 -14191
rect -3429 -14198 -161 -14195
rect 161 -14198 3429 -14195
rect -3429 -14233 3429 -14198
rect -3252 -14272 3252 -14233
rect -3075 -14309 3075 -14272
rect -2898 -14344 2898 -14309
rect -2720 -14377 2720 -14344
rect -2541 -14408 2541 -14377
rect -2363 -14436 2363 -14408
rect -2184 -14462 2184 -14436
rect -2004 -14486 2004 -14462
rect -1825 -14508 1825 -14486
rect -1645 -14527 1645 -14508
rect -1465 -14544 1465 -14527
rect -1284 -14559 1284 -14544
rect -1104 -14571 1104 -14559
rect -923 -14581 923 -14571
rect -742 -14589 742 -14581
rect -561 -14595 561 -14589
rect -380 -14598 380 -14595
rect -200 -14600 199 -14598
use skullfet_inverter_5v  skullfet_inverter_0
timestamp 1735296207
transform 1 0 11000 0 1 -1400
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_1
timestamp 1735296207
transform -1 0 12466 0 1 2136
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_2
timestamp 1735296207
transform 1 0 8914 0 1 5358
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_3
timestamp 1735296207
transform 1 0 6480 0 1 7980
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_4
timestamp 1735296207
transform 1 0 3384 0 1 9770
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_5
timestamp 1735296207
transform 1 0 -104 0 1 10566
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_6
timestamp 1735296207
transform 1 0 -3670 0 1 10298
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_7
timestamp 1735296207
transform 1 0 -6998 0 1 8992
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_8
timestamp 1735296207
transform 1 0 -9796 0 1 6762
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_9
timestamp 1735296207
transform 1 0 -11810 0 1 3806
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_10
timestamp 1735296207
transform -1 0 -10864 0 1 388
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_11
timestamp 1735296207
transform 1 0 -12864 0 1 -3188
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_12
timestamp 1735296207
transform -1 0 -9810 0 1 -6606
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_13
timestamp 1735296207
transform -1 0 -7796 0 -1 -6762
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_14
timestamp 1735296207
transform -1 0 -5000 0 -1 -8992
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_15
timestamp 1735296207
transform -1 0 -1670 0 -1 -10298
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_16
timestamp 1735296207
transform -1 0 1896 0 -1 -10566
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_17
timestamp 1735296207
transform -1 0 5384 0 -1 -9770
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_18
timestamp 1735296207
transform -1 0 8480 0 -1 -7980
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_19
timestamp 1735296207
transform -1 0 10914 0 1 -8158
box 454 132 2110 3088
use skullfet_inverter_5v  skullfet_inverter_20
timestamp 1735296207
transform -1 0 12466 0 1 -4936
box 454 132 2110 3088
<< end >>
