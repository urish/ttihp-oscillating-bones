* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7] VDPWR VGND
X0 a_13289_43697# uo_out[2].t2 VDPWR.t37 VDPWR.t36 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_16868_43697# a_17160_43997# a_17111_44089# VDPWR.t85 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2 a_16596_43697# a_16868_43697# VGND.t66 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VDPWR.t101 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VDPWR.t100 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X4 VGND.t20 uo_out[0].t2 ring_0/skullfet_inverter_6.A VGND.t19 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X5 VGND.t30 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X6 VGND.t80 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t79 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X7 a_15221_43697# uo_out[1].t2 VDPWR.t23 VDPWR.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X8 VDPWR.t61 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VDPWR.t60 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X9 a_15179_44089# a_14664_43697# VDPWR.t35 VDPWR.t34 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X10 a_17360_43697# a_17160_43997# a_17509_43723# VGND.t63 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X11 VGND.t57 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VGND.t56 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X12 ring_0/skullfet_inverter_6.A uo_out[0].t3 VDPWR.t27 VDPWR.t26 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X13 a_15577_43723# a_15357_43723# VGND.t78 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X14 VGND.t28 a_14664_43697# uo_out[2].t0 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VDPWR.t55 a_13289_43697# a_13296_43997# VDPWR.t54 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 VGND.t60 a_15221_43697# a_15228_43997# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t77 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t76 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X18 a_13843_43723# a_13296_43997# a_13496_43697# VDPWR.t69 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X19 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VDPWR.t109 VDPWR.t108 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X20 VGND.t10 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_8.A VGND.t9 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X21 a_16501_43697# a_16596_43697# VGND.t34 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X22 a_12637_43697# a_12732_43697# VDPWR.t5 VDPWR.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X23 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t18 VGND.t17 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X24 VGND.t62 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t61 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X25 a_17289_43723# a_17153_43697# a_16868_43697# VDPWR.t89 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 a_13224_43723# a_12732_43697# VGND.t5 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VDPWR.t33 a_14664_43697# uo_out[2].t1 VDPWR.t32 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t45 VGND.t44 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X29 VDPWR.t49 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VDPWR.t48 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X30 VGND.t71 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t70 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X31 VGND.t73 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t72 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X32 a_15156_43723# a_14664_43697# VGND.t27 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X33 a_17707_43723# a_17153_43697# a_17360_43697# VGND.t65 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X34 a_14936_43697# a_15228_43997# a_15179_44089# VDPWR.t67 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X35 a_13289_43697# uo_out[2].t3 VGND.t29 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X36 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_7.A VDPWR.t11 VDPWR.t10 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X37 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VDPWR.t83 VDPWR.t82 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X38 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VDPWR.t97 VDPWR.t96 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X39 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_8.A VDPWR.t9 VDPWR.t8 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X40 VGND.t43 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X41 a_14664_43697# a_14936_43697# VGND.t82 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X42 VGND.t74 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X43 VGND.t12 a_13496_43697# a_13425_43723# VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X44 a_13247_44089# a_12732_43697# VDPWR.t3 VDPWR.t2 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X45 a_15221_43697# uo_out[1].t3 VGND.t23 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X46 a_15428_43697# a_15228_43997# a_15577_43723# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X47 a_13645_43723# a_13425_43723# VGND.t39 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X48 VDPWR.t17 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VDPWR.t16 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X49 VDPWR.t47 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VDPWR.t46 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X50 VGND.t81 a_15428_43697# a_15357_43723# VGND.t11 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X51 VGND.t3 a_12732_43697# uo_out[3].t0 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X52 VGND.t68 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t67 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X53 VDPWR.t77 a_17360_43697# a_17289_43723# VDPWR.t76 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X54 a_16868_43697# a_17153_43697# a_17088_43723# VGND.t63 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X55 a_14664_43697# a_14936_43697# VDPWR.t113 VDPWR.t112 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X56 VGND.t41 a_13289_43697# a_13296_43997# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X57 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VDPWR.t99 VDPWR.t98 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X58 VDPWR.t19 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VDPWR.t18 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X59 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VDPWR.t75 VDPWR.t74 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X60 a_14569_43697# a_14664_43697# VGND.t26 VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X61 a_15604_44089# a_15357_43723# VDPWR.t107 VDPWR.t106 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X62 a_15357_43723# a_15221_43697# a_14936_43697# VDPWR.t81 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X63 a_15428_43697# a_15221_43697# a_15604_44089# VDPWR.t80 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X64 a_12732_43697# a_13004_43697# VGND.t69 VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X65 VGND.t49 ring_0/skullfet_inverter_4.A uo_out[0].t0 VGND.t48 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X66 VDPWR.t57 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VDPWR.t56 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X67 VDPWR.t1 a_12732_43697# uo_out[3].t1 VDPWR.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X68 VGND.t22 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t21 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X69 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VDPWR.t65 VDPWR.t64 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X70 VDPWR.t71 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VDPWR.t70 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X71 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VDPWR.t93 VDPWR.t92 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X72 a_17289_43723# a_17160_43997# a_16868_43697# VGND.t63 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X73 a_17153_43697# uo_out[0].t4 VDPWR.t25 VDPWR.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X74 a_17536_44089# a_17289_43723# VDPWR.t29 VDPWR.t28 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X75 a_17360_43697# a_17153_43697# a_17536_44089# VDPWR.t88 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X76 a_17111_44089# a_16596_43697# VDPWR.t45 VDPWR.t44 sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X77 a_15775_43723# a_15221_43697# a_15428_43697# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X78 a_13004_43697# a_13296_43997# a_13247_44089# VDPWR.t68 sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X79 VDPWR.t7 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VDPWR.t6 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X80 a_12732_43697# a_13004_43697# VDPWR.t95 VDPWR.t94 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X81 VGND.t14 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t13 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X82 VGND.t75 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X83 uo_out[0].t1 ring_0/skullfet_inverter_4.A VDPWR.t63 VDPWR.t62 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X84 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VDPWR.t21 VDPWR.t20 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X85 a_16501_43697# a_16596_43697# VDPWR.t43 VDPWR.t42 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X86 a_13496_43697# a_13296_43997# a_13645_43723# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X87 VDPWR.t87 a_17153_43697# a_17160_43997# VDPWR.t86 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X88 VDPWR.t111 a_15428_43697# a_15357_43723# VDPWR.t110 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X89 VGND.t51 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t50 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X90 a_14936_43697# a_15221_43697# a_15156_43723# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X91 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VDPWR.t15 VDPWR.t14 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X92 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t53 VGND.t52 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X93 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VDPWR.t73 VDPWR.t72 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X94 a_12637_43697# a_12732_43697# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X95 a_13672_44089# a_13425_43723# VDPWR.t51 VDPWR.t50 sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X96 a_13425_43723# a_13296_43997# a_13004_43697# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X97 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X98 a_13425_43723# a_13289_43697# a_13004_43697# VDPWR.t53 sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 a_13496_43697# a_13289_43697# a_13672_44089# VDPWR.t52 sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X100 VDPWR.t39 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VDPWR.t38 sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X101 VDPWR.t103 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VDPWR.t102 sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X102 VDPWR.t59 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VDPWR.t58 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X103 a_15357_43723# a_15228_43997# a_14936_43697# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X104 a_17153_43697# uo_out[0].t5 VGND.t46 VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X105 a_17509_43723# a_17289_43723# VGND.t25 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X106 VGND.t33 a_16596_43697# uo_out[1].t0 VGND.t32 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X107 a_13843_43723# a_13289_43697# a_13496_43697# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X108 VGND.t59 a_17360_43697# a_17289_43723# VGND.t58 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X109 VGND.t6 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t2 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X110 VDPWR.t79 a_15221_43697# a_15228_43997# VDPWR.t78 sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X111 VGND.t47 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VGND.t4 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X112 a_15775_43723# a_15228_43997# a_15428_43697# VDPWR.t66 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X113 a_13004_43697# a_13289_43697# a_13224_43723# VGND.t40 sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X114 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t36 VGND.t35 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X115 a_16596_43697# a_16868_43697# VDPWR.t91 VDPWR.t90 sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X116 a_14569_43697# a_14664_43697# VDPWR.t31 VDPWR.t30 sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X117 VGND.t55 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VGND.t54 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X118 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t16 VGND.t15 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X119 a_17707_43723# a_17160_43997# a_17360_43697# VDPWR.t84 sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X120 VDPWR.t41 a_16596_43697# uo_out[1].t1 VDPWR.t40 sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X121 VGND.t8 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_9.A VGND.t7 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X122 VDPWR.t13 a_13496_43697# a_13425_43723# VDPWR.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X123 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VDPWR.t105 VDPWR.t104 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X124 VGND.t64 a_17153_43697# a_17160_43997# VGND.t42 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X125 a_17088_43723# a_16596_43697# VGND.t31 VGND.t24 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 uo_out[2].n2 uo_out[2].t1 313.104
R1 uo_out[2].n0 uo_out[2].t2 294.557
R2 uo_out[2].t0 uo_out[2].n2 265.769
R3 uo_out[2] uo_out[2].t0 262.318
R4 uo_out[2].n0 uo_out[2].t3 211.01
R5 uo_out[2].n1 uo_out[2].n0 152
R6 uo_out[2].n5 uo_out[2] 16.2155
R7 uo_out[2].n4 uo_out[2].n1 11.6311
R8 uo_out[2].n4 uo_out[2].n3 9.3005
R9 uo_out[2].n3 uo_out[2] 7.17626
R10 uo_out[2].n3 uo_out[2].n2 4.84898
R11 uo_out[2].n5 uo_out[2].n4 4.51042
R12 uo_out[2].n1 uo_out[2] 1.37896
R13 uo_out[2] uo_out[2].n5 0.0730806
R14 VDPWR.n5 VDPWR.t109 739.681
R15 VDPWR.n3 VDPWR.t71 739.681
R16 VDPWR.n230 VDPWR.t17 739.681
R17 VDPWR.n227 VDPWR.t73 739.681
R18 VDPWR.n224 VDPWR.t97 739.681
R19 VDPWR.n366 VDPWR.t21 739.681
R20 VDPWR.n278 VDPWR.t47 739.681
R21 VDPWR.n280 VDPWR.t75 739.681
R22 VDPWR.n228 VDPWR.t49 739.681
R23 VDPWR.n232 VDPWR.t19 739.681
R24 VDPWR.n0 VDPWR.t59 739.681
R25 VDPWR.n7 VDPWR.t83 739.681
R26 VDPWR.n225 VDPWR.t99 739.681
R27 VDPWR.n222 VDPWR.t105 739.681
R28 VDPWR.n177 VDPWR.t27 739.681
R29 VDPWR.n173 VDPWR.t93 739.681
R30 VDPWR.n152 VDPWR.t11 739.681
R31 VDPWR.n360 VDPWR.t9 739.681
R32 VDPWR.n363 VDPWR.t65 739.681
R33 VDPWR.n199 VDPWR.t63 739.681
R34 VDPWR.n288 VDPWR.t15 739.681
R35 VDPWR.n7 VDPWR.t82 707.852
R36 VDPWR.n5 VDPWR.t108 707.852
R37 VDPWR.n3 VDPWR.t70 707.852
R38 VDPWR.n230 VDPWR.t16 707.852
R39 VDPWR.n227 VDPWR.t72 707.852
R40 VDPWR.n225 VDPWR.t98 707.852
R41 VDPWR.n224 VDPWR.t96 707.852
R42 VDPWR.n222 VDPWR.t104 707.852
R43 VDPWR.n177 VDPWR.t26 707.852
R44 VDPWR.n173 VDPWR.t92 707.852
R45 VDPWR.n152 VDPWR.t10 707.852
R46 VDPWR.n360 VDPWR.t8 707.852
R47 VDPWR.n363 VDPWR.t64 707.852
R48 VDPWR.n366 VDPWR.t20 707.852
R49 VDPWR.n199 VDPWR.t62 707.852
R50 VDPWR.n288 VDPWR.t14 707.852
R51 VDPWR.n278 VDPWR.t46 707.852
R52 VDPWR.n280 VDPWR.t74 707.852
R53 VDPWR.n228 VDPWR.t48 707.852
R54 VDPWR.n232 VDPWR.t18 707.852
R55 VDPWR.n0 VDPWR.t58 707.852
R56 VDPWR.n92 VDPWR.t3 667.734
R57 VDPWR.n60 VDPWR.t35 667.734
R58 VDPWR.n130 VDPWR.t45 667.734
R59 VDPWR.n107 VDPWR.t61 666.677
R60 VDPWR.n46 VDPWR.t103 666.677
R61 VDPWR.n144 VDPWR.t57 666.677
R62 VDPWR.t90 VDPWR.t44 624.456
R63 VDPWR.t34 VDPWR.t112 624.456
R64 VDPWR.t2 VDPWR.t94 624.456
R65 VDPWR.n110 VDPWR.n109 604.394
R66 VDPWR.n39 VDPWR.n38 604.394
R67 VDPWR.n148 VDPWR.n10 604.394
R68 VDPWR.t56 VDPWR.t86 556.386
R69 VDPWR.t42 VDPWR.t40 556.386
R70 VDPWR.t78 VDPWR.t102 556.386
R71 VDPWR.t32 VDPWR.t30 556.386
R72 VDPWR.t54 VDPWR.t60 556.386
R73 VDPWR.t0 VDPWR.t4 556.386
R74 VDPWR.n118 VDPWR.t6 414.33
R75 VDPWR.t38 VDPWR.n116 414.33
R76 VDPWR.t76 VDPWR.t28 390.654
R77 VDPWR.t106 VDPWR.t110 390.654
R78 VDPWR.t50 VDPWR.t12 390.654
R79 VDPWR.t44 VDPWR.t85 337.384
R80 VDPWR.t67 VDPWR.t34 337.384
R81 VDPWR.t68 VDPWR.t2 337.384
R82 VDPWR.n90 VDPWR.n80 333.348
R83 VDPWR.n62 VDPWR.n30 333.348
R84 VDPWR.n18 VDPWR.n17 333.348
R85 VDPWR.n76 VDPWR.n75 320.976
R86 VDPWR.n53 VDPWR.n34 320.976
R87 VDPWR.n137 VDPWR.n14 320.976
R88 VDPWR.t28 VDPWR.t88 304.829
R89 VDPWR.t80 VDPWR.t106 304.829
R90 VDPWR.t52 VDPWR.t50 304.829
R91 VDPWR.t6 VDPWR.t42 287.072
R92 VDPWR.t30 VDPWR.t38 287.072
R93 VDPWR.t4 VDPWR.t100 287.072
R94 VDPWR.t88 VDPWR.t84 281.154
R95 VDPWR.t89 VDPWR.t76 281.154
R96 VDPWR.t66 VDPWR.t80 281.154
R97 VDPWR.t110 VDPWR.t81 281.154
R98 VDPWR.t69 VDPWR.t52 281.154
R99 VDPWR.t12 VDPWR.t53 281.154
R100 VDPWR.n118 VDPWR.n117 272.274
R101 VDPWR.n117 VDPWR 272.274
R102 VDPWR.n116 VDPWR.n115 272.274
R103 VDPWR.n115 VDPWR 272.274
R104 VDPWR.t84 VDPWR.t56 251.559
R105 VDPWR.t102 VDPWR.t66 251.559
R106 VDPWR.t60 VDPWR.t69 251.559
R107 VDPWR.t86 VDPWR.t24 248.599
R108 VDPWR.t85 VDPWR.t89 248.599
R109 VDPWR.t40 VDPWR.t90 248.599
R110 VDPWR.t22 VDPWR.t78 248.599
R111 VDPWR.t81 VDPWR.t67 248.599
R112 VDPWR.t112 VDPWR.t32 248.599
R113 VDPWR.t36 VDPWR.t54 248.599
R114 VDPWR.t53 VDPWR.t68 248.599
R115 VDPWR.t94 VDPWR.t0 248.599
R116 VDPWR.n84 VDPWR.n83 240.522
R117 VDPWR.n68 VDPWR.n27 240.522
R118 VDPWR.n21 VDPWR.n20 240.522
R119 VDPWR.n115 VDPWR.n114 213.119
R120 VDPWR.n116 VDPWR.n24 213.119
R121 VDPWR.n117 VDPWR.n22 213.119
R122 VDPWR.n119 VDPWR.n118 213.119
R123 VDPWR.n75 VDPWR.t51 113.98
R124 VDPWR.n34 VDPWR.t107 113.98
R125 VDPWR.n14 VDPWR.t29 113.98
R126 VDPWR.t24 VDPWR 91.745
R127 VDPWR VDPWR.t22 91.745
R128 VDPWR VDPWR.t36 91.745
R129 VDPWR.n83 VDPWR.t5 61.9872
R130 VDPWR.n27 VDPWR.t31 61.9872
R131 VDPWR.n20 VDPWR.t43 61.9872
R132 VDPWR.n109 VDPWR.t37 41.5552
R133 VDPWR.n109 VDPWR.t55 41.5552
R134 VDPWR.n38 VDPWR.t23 41.5552
R135 VDPWR.n38 VDPWR.t79 41.5552
R136 VDPWR.n10 VDPWR.t25 41.5552
R137 VDPWR.n10 VDPWR.t87 41.5552
R138 VDPWR.n75 VDPWR.t13 35.4605
R139 VDPWR.n34 VDPWR.t111 35.4605
R140 VDPWR.n14 VDPWR.t77 35.4605
R141 VDPWR.n89 VDPWR.n81 34.6358
R142 VDPWR.n85 VDPWR.n81 34.6358
R143 VDPWR.n103 VDPWR.n73 34.6358
R144 VDPWR.n103 VDPWR.n102 34.6358
R145 VDPWR.n102 VDPWR.n101 34.6358
R146 VDPWR.n98 VDPWR.n97 34.6358
R147 VDPWR.n97 VDPWR.n96 34.6358
R148 VDPWR.n96 VDPWR.n78 34.6358
R149 VDPWR.n63 VDPWR.n28 34.6358
R150 VDPWR.n67 VDPWR.n28 34.6358
R151 VDPWR.n48 VDPWR.n47 34.6358
R152 VDPWR.n48 VDPWR.n35 34.6358
R153 VDPWR.n52 VDPWR.n35 34.6358
R154 VDPWR.n55 VDPWR.n54 34.6358
R155 VDPWR.n55 VDPWR.n32 34.6358
R156 VDPWR.n59 VDPWR.n32 34.6358
R157 VDPWR.n126 VDPWR.n125 34.6358
R158 VDPWR.n125 VDPWR.n124 34.6358
R159 VDPWR.n143 VDPWR.n142 34.6358
R160 VDPWR.n142 VDPWR.n12 34.6358
R161 VDPWR.n138 VDPWR.n12 34.6358
R162 VDPWR.n136 VDPWR.n135 34.6358
R163 VDPWR.n135 VDPWR.n15 34.6358
R164 VDPWR.n131 VDPWR.n15 34.6358
R165 VDPWR.n91 VDPWR.n90 32.0005
R166 VDPWR.n62 VDPWR.n61 32.0005
R167 VDPWR.n129 VDPWR.n18 32.0005
R168 VDPWR.n149 VDPWR.n148 30.7593
R169 VDPWR.n92 VDPWR.n91 30.4946
R170 VDPWR.n61 VDPWR.n60 30.4946
R171 VDPWR.n130 VDPWR.n129 30.4946
R172 VDPWR.n83 VDPWR.t101 30.1692
R173 VDPWR.n27 VDPWR.t39 30.1692
R174 VDPWR.n20 VDPWR.t7 30.1692
R175 VDPWR.n107 VDPWR.n73 27.4829
R176 VDPWR.n69 VDPWR.n68 27.4829
R177 VDPWR.n47 VDPWR.n46 27.4829
R178 VDPWR.n120 VDPWR.n21 27.4829
R179 VDPWR.n144 VDPWR.n143 27.4829
R180 VDPWR.n80 VDPWR.t95 26.5955
R181 VDPWR.n80 VDPWR.t1 26.5955
R182 VDPWR.n30 VDPWR.t113 26.5955
R183 VDPWR.n30 VDPWR.t33 26.5955
R184 VDPWR.n17 VDPWR.t91 26.5955
R185 VDPWR.n17 VDPWR.t41 26.5955
R186 VDPWR.n85 VDPWR.n84 25.6005
R187 VDPWR.n68 VDPWR.n67 25.6005
R188 VDPWR.n124 VDPWR.n21 25.6005
R189 VDPWR.n114 VDPWR.n25 23.7181
R190 VDPWR.n69 VDPWR.n24 23.7181
R191 VDPWR.n41 VDPWR.n22 23.7181
R192 VDPWR.n120 VDPWR.n119 23.7181
R193 VDPWR.n110 VDPWR.n108 22.9652
R194 VDPWR.n45 VDPWR.n39 22.9652
R195 VDPWR.n148 VDPWR.n9 22.9652
R196 VDPWR.n108 VDPWR.n107 21.8358
R197 VDPWR.n46 VDPWR.n45 21.8358
R198 VDPWR.n144 VDPWR.n9 21.8358
R199 VDPWR.n110 VDPWR.n25 21.4593
R200 VDPWR.n41 VDPWR.n39 21.4593
R201 VDPWR.n101 VDPWR.n76 18.4476
R202 VDPWR.n53 VDPWR.n52 18.4476
R203 VDPWR.n138 VDPWR.n137 18.4476
R204 VDPWR.n150 VDPWR.n149 16.5693
R205 VDPWR.n98 VDPWR.n76 16.1887
R206 VDPWR.n54 VDPWR.n53 16.1887
R207 VDPWR.n137 VDPWR.n136 16.1887
R208 VDPWR.n92 VDPWR.n78 15.0593
R209 VDPWR.n60 VDPWR.n59 15.0593
R210 VDPWR.n131 VDPWR.n130 15.0593
R211 VDPWR.n8 VDPWR.n7 13.377
R212 VDPWR.n226 VDPWR.n225 13.377
R213 VDPWR.n223 VDPWR.n222 13.377
R214 VDPWR.n178 VDPWR.n177 13.377
R215 VDPWR.n174 VDPWR.n173 13.377
R216 VDPWR.n153 VDPWR.n152 13.377
R217 VDPWR.n361 VDPWR.n360 13.377
R218 VDPWR.n364 VDPWR.n363 13.377
R219 VDPWR.n200 VDPWR.n199 13.377
R220 VDPWR.n289 VDPWR.n288 13.377
R221 VDPWR VDPWR.n5 13.3202
R222 VDPWR.n4 VDPWR.n3 13.3202
R223 VDPWR.n231 VDPWR.n230 13.3202
R224 VDPWR VDPWR.n227 13.3202
R225 VDPWR VDPWR.n224 13.3202
R226 VDPWR VDPWR.n366 13.3202
R227 VDPWR.n279 VDPWR.n278 13.3202
R228 VDPWR VDPWR.n280 13.3202
R229 VDPWR.n229 VDPWR.n228 13.3202
R230 VDPWR.n233 VDPWR.n232 13.3202
R231 VDPWR.n373 VDPWR.n0 13.3202
R232 VDPWR.n114 VDPWR.n24 12.8005
R233 VDPWR.n119 VDPWR.n22 12.8005
R234 VDPWR.n283 VDPWR 9.7375
R235 VDPWR.n281 VDPWR 9.39357
R236 VDPWR.n148 VDPWR.n147 9.3005
R237 VDPWR.n146 VDPWR.n9 9.3005
R238 VDPWR.n145 VDPWR.n144 9.3005
R239 VDPWR.n143 VDPWR.n11 9.3005
R240 VDPWR.n142 VDPWR.n141 9.3005
R241 VDPWR.n140 VDPWR.n12 9.3005
R242 VDPWR.n139 VDPWR.n138 9.3005
R243 VDPWR.n136 VDPWR.n13 9.3005
R244 VDPWR.n135 VDPWR.n134 9.3005
R245 VDPWR.n133 VDPWR.n15 9.3005
R246 VDPWR.n132 VDPWR.n131 9.3005
R247 VDPWR.n130 VDPWR.n16 9.3005
R248 VDPWR.n129 VDPWR.n128 9.3005
R249 VDPWR.n127 VDPWR.n126 9.3005
R250 VDPWR.n125 VDPWR.n19 9.3005
R251 VDPWR.n124 VDPWR.n123 9.3005
R252 VDPWR.n122 VDPWR.n21 9.3005
R253 VDPWR.n121 VDPWR.n120 9.3005
R254 VDPWR.n119 VDPWR.n23 9.3005
R255 VDPWR.n40 VDPWR.n22 9.3005
R256 VDPWR.n42 VDPWR.n41 9.3005
R257 VDPWR.n43 VDPWR.n39 9.3005
R258 VDPWR.n45 VDPWR.n44 9.3005
R259 VDPWR.n46 VDPWR.n37 9.3005
R260 VDPWR.n47 VDPWR.n36 9.3005
R261 VDPWR.n49 VDPWR.n48 9.3005
R262 VDPWR.n50 VDPWR.n35 9.3005
R263 VDPWR.n52 VDPWR.n51 9.3005
R264 VDPWR.n54 VDPWR.n33 9.3005
R265 VDPWR.n56 VDPWR.n55 9.3005
R266 VDPWR.n57 VDPWR.n32 9.3005
R267 VDPWR.n59 VDPWR.n58 9.3005
R268 VDPWR.n60 VDPWR.n31 9.3005
R269 VDPWR.n61 VDPWR.n29 9.3005
R270 VDPWR.n64 VDPWR.n63 9.3005
R271 VDPWR.n65 VDPWR.n28 9.3005
R272 VDPWR.n67 VDPWR.n66 9.3005
R273 VDPWR.n68 VDPWR.n26 9.3005
R274 VDPWR.n70 VDPWR.n69 9.3005
R275 VDPWR.n71 VDPWR.n24 9.3005
R276 VDPWR.n114 VDPWR.n113 9.3005
R277 VDPWR.n112 VDPWR.n25 9.3005
R278 VDPWR.n111 VDPWR.n110 9.3005
R279 VDPWR.n108 VDPWR.n72 9.3005
R280 VDPWR.n107 VDPWR.n106 9.3005
R281 VDPWR.n105 VDPWR.n73 9.3005
R282 VDPWR.n104 VDPWR.n103 9.3005
R283 VDPWR.n102 VDPWR.n74 9.3005
R284 VDPWR.n101 VDPWR.n100 9.3005
R285 VDPWR.n99 VDPWR.n98 9.3005
R286 VDPWR.n97 VDPWR.n77 9.3005
R287 VDPWR.n96 VDPWR.n95 9.3005
R288 VDPWR.n94 VDPWR.n78 9.3005
R289 VDPWR.n93 VDPWR.n92 9.3005
R290 VDPWR.n91 VDPWR.n79 9.3005
R291 VDPWR.n89 VDPWR.n88 9.3005
R292 VDPWR.n87 VDPWR.n81 9.3005
R293 VDPWR.n86 VDPWR.n85 9.3005
R294 VDPWR.n369 VDPWR.n8 8.51977
R295 VDPWR.n285 VDPWR 8.13646
R296 VDPWR.n282 VDPWR.n277 7.53241
R297 VDPWR.n365 VDPWR.n364 7.53109
R298 VDPWR.n362 VDPWR.n361 7.45619
R299 VDPWR.n84 VDPWR.n82 7.4049
R300 VDPWR.n6 VDPWR 7.19357
R301 VDPWR.n358 VDPWR.n153 6.79323
R302 VDPWR.n284 VDPWR.n226 6.76538
R303 VDPWR.n367 VDPWR 6.40107
R304 VDPWR.n277 VDPWR.n229 6.34337
R305 VDPWR.n276 VDPWR.n231 6.19552
R306 VDPWR.n281 VDPWR.n279 6.1805
R307 VDPWR.n286 VDPWR.n223 6.08268
R308 VDPWR.n283 VDPWR.n282 6.07848
R309 VDPWR.n175 VDPWR.n174 6.01772
R310 VDPWR.n290 VDPWR.n289 6.01019
R311 VDPWR.n312 VDPWR.n200 5.71852
R312 VDPWR.n333 VDPWR.n178 5.65925
R313 VDPWR.n234 VDPWR.n233 5.44488
R314 VDPWR.n373 VDPWR.n372 5.3655
R315 VDPWR.n6 VDPWR.n4 5.233
R316 VDPWR.n287 VDPWR.n286 4.1734
R317 VDPWR.n370 VDPWR.n369 4.09754
R318 VDPWR.n150 VDPWR 3.44278
R319 VDPWR.n334 VDPWR.n176 3.07281
R320 VDPWR.n90 VDPWR.n89 2.63579
R321 VDPWR.n63 VDPWR.n62 2.63579
R322 VDPWR.n126 VDPWR.n18 2.63579
R323 VDPWR.n368 VDPWR.n150 1.94486
R324 VDPWR.n282 VDPWR.n281 1.25038
R325 VDPWR.n371 VDPWR.n370 1.04464
R326 VDPWR.n277 VDPWR.n276 0.897709
R327 VDPWR.n367 VDPWR.n365 0.877511
R328 VDPWR.n218 VDPWR.n217 0.861295
R329 VDPWR.n369 VDPWR.n368 0.848036
R330 VDPWR.n286 VDPWR.n285 0.838747
R331 VDPWR.n284 VDPWR.n283 0.83329
R332 VDPWR.n285 VDPWR.n284 0.810795
R333 VDPWR.n362 VDPWR.n359 0.698295
R334 VDPWR.n276 VDPWR.n275 0.574375
R335 VDPWR.n365 VDPWR.n362 0.53699
R336 VDPWR.n219 VDPWR.n218 0.507602
R337 VDPWR.n335 VDPWR.n334 0.491158
R338 VDPWR.n370 VDPWR.n6 0.456575
R339 VDPWR.n220 VDPWR.n219 0.391496
R340 VDPWR.n179 VDPWR.n176 0.380996
R341 VDPWR.n221 VDPWR.n220 0.325974
R342 VDPWR.n275 VDPWR.n234 0.323617
R343 VDPWR.n287 VDPWR.n221 0.320751
R344 VDPWR.n180 VDPWR.n179 0.263105
R345 VDPWR.n181 VDPWR.n180 0.23221
R346 VDPWR.n291 VDPWR.n221 0.198913
R347 VDPWR.n292 VDPWR.n220 0.195812
R348 VDPWR.n182 VDPWR.n181 0.193814
R349 VDPWR.n293 VDPWR.n219 0.192808
R350 VDPWR.n294 VDPWR.n218 0.189894
R351 VDPWR.n183 VDPWR.n182 0.183989
R352 VDPWR.n359 VDPWR.n151 0.169675
R353 VDPWR.n336 VDPWR.n335 0.168706
R354 VDPWR.n332 VDPWR.n176 0.162658
R355 VDPWR.n184 VDPWR.n183 0.157627
R356 VDPWR.n82 VDPWR 0.156264
R357 VDPWR.n358 VDPWR.n357 0.154418
R358 VDPWR.n296 VDPWR.n295 0.154418
R359 VDPWR.n310 VDPWR.n202 0.153485
R360 VDPWR.n185 VDPWR.n184 0.148565
R361 VDPWR.n254 VDPWR.n1 0.147626
R362 VDPWR.n86 VDPWR.n82 0.144904
R363 VDPWR.n331 VDPWR.n179 0.143882
R364 VDPWR.n330 VDPWR.n180 0.142412
R365 VDPWR.n328 VDPWR.n182 0.140206
R366 VDPWR.n329 VDPWR.n181 0.140035
R367 VDPWR.n326 VDPWR.n184 0.139637
R368 VDPWR.n327 VDPWR.n183 0.139471
R369 VDPWR.n272 VDPWR.n235 0.137548
R370 VDPWR.n324 VDPWR.n186 0.137405
R371 VDPWR.n325 VDPWR.n185 0.137265
R372 VDPWR.n270 VDPWR.n237 0.136933
R373 VDPWR.n323 VDPWR.n187 0.136661
R374 VDPWR.n274 VDPWR.n273 0.136661
R375 VDPWR.n356 VDPWR.n355 0.136529
R376 VDPWR.n297 VDPWR.n215 0.136529
R377 VDPWR.n271 VDPWR.n236 0.136042
R378 VDPWR.n322 VDPWR.n188 0.135917
R379 VDPWR.n186 VDPWR.n185 0.135794
R380 VDPWR.n337 VDPWR.n171 0.135785
R381 VDPWR.n255 VDPWR.n252 0.135774
R382 VDPWR.n266 VDPWR.n241 0.135656
R383 VDPWR.n357 VDPWR.n151 0.13561
R384 VDPWR.n296 VDPWR.n216 0.13561
R385 VDPWR.n267 VDPWR.n240 0.135531
R386 VDPWR.n269 VDPWR.n238 0.135409
R387 VDPWR.n259 VDPWR.n248 0.135368
R388 VDPWR.n353 VDPWR.n155 0.135321
R389 VDPWR.n299 VDPWR.n213 0.135321
R390 VDPWR.n320 VDPWR.n190 0.135289
R391 VDPWR.n261 VDPWR.n246 0.13524
R392 VDPWR.n264 VDPWR.n243 0.134994
R393 VDPWR.n254 VDPWR.n253 0.134918
R394 VDPWR.n257 VDPWR.n250 0.134667
R395 VDPWR.n321 VDPWR.n189 0.134429
R396 VDPWR.n263 VDPWR.n244 0.134203
R397 VDPWR.n318 VDPWR.n192 0.133884
R398 VDPWR.n317 VDPWR.n193 0.133884
R399 VDPWR.n268 VDPWR.n239 0.133884
R400 VDPWR.n319 VDPWR.n191 0.133783
R401 VDPWR.n343 VDPWR.n165 0.133617
R402 VDPWR.n309 VDPWR.n203 0.133617
R403 VDPWR.n354 VDPWR.n154 0.133536
R404 VDPWR.n298 VDPWR.n214 0.133536
R405 VDPWR.n351 VDPWR.n157 0.133312
R406 VDPWR.n338 VDPWR.n170 0.133312
R407 VDPWR.n314 VDPWR.n196 0.133312
R408 VDPWR.n301 VDPWR.n211 0.133312
R409 VDPWR.n303 VDPWR.n209 0.133205
R410 VDPWR.n348 VDPWR.n160 0.133101
R411 VDPWR.n256 VDPWR.n251 0.133
R412 VDPWR.n345 VDPWR.n163 0.132901
R413 VDPWR.n307 VDPWR.n205 0.132901
R414 VDPWR.n258 VDPWR.n249 0.132901
R415 VDPWR.n340 VDPWR.n168 0.13262
R416 VDPWR.n312 VDPWR.n198 0.13262
R417 VDPWR.n262 VDPWR.n245 0.13262
R418 VDPWR.n315 VDPWR.n195 0.132444
R419 VDPWR.n265 VDPWR.n242 0.132444
R420 VDPWR.n316 VDPWR.n194 0.13236
R421 VDPWR.n350 VDPWR.n158 0.132349
R422 VDPWR.n302 VDPWR.n210 0.132349
R423 VDPWR.n347 VDPWR.n161 0.132167
R424 VDPWR.n305 VDPWR.n207 0.132167
R425 VDPWR.n260 VDPWR.n247 0.13191
R426 VDPWR.n341 VDPWR.n167 0.131829
R427 VDPWR.n273 VDPWR.n272 0.131701
R428 VDPWR.n352 VDPWR.n156 0.131576
R429 VDPWR.n300 VDPWR.n212 0.131576
R430 VDPWR.n349 VDPWR.n159 0.131412
R431 VDPWR.n304 VDPWR.n208 0.131333
R432 VDPWR.n346 VDPWR.n162 0.131257
R433 VDPWR.n306 VDPWR.n206 0.131257
R434 VDPWR.n339 VDPWR.n169 0.130901
R435 VDPWR.n313 VDPWR.n197 0.130901
R436 VDPWR.n371 VDPWR.n2 0.130781
R437 VDPWR.n342 VDPWR.n166 0.130247
R438 VDPWR.n272 VDPWR.n271 0.130144
R439 VDPWR.n187 VDPWR.n186 0.130052
R440 VDPWR.n344 VDPWR.n164 0.129506
R441 VDPWR.n308 VDPWR.n204 0.129506
R442 VDPWR.n336 VDPWR.n172 0.12922
R443 VDPWR.n355 VDPWR.n151 0.124945
R444 VDPWR.n216 VDPWR.n215 0.124945
R445 VDPWR.n188 VDPWR.n187 0.12426
R446 VDPWR.n355 VDPWR.n354 0.122959
R447 VDPWR.n215 VDPWR.n214 0.122959
R448 VDPWR.n271 VDPWR.n270 0.122756
R449 VDPWR.n270 VDPWR.n269 0.122197
R450 VDPWR.n202 VDPWR.n201 0.121074
R451 VDPWR.n147 VDPWR.n146 0.120292
R452 VDPWR.n146 VDPWR.n145 0.120292
R453 VDPWR.n145 VDPWR.n11 0.120292
R454 VDPWR.n141 VDPWR.n11 0.120292
R455 VDPWR.n141 VDPWR.n140 0.120292
R456 VDPWR.n140 VDPWR.n139 0.120292
R457 VDPWR.n139 VDPWR.n13 0.120292
R458 VDPWR.n134 VDPWR.n13 0.120292
R459 VDPWR.n134 VDPWR.n133 0.120292
R460 VDPWR.n133 VDPWR.n132 0.120292
R461 VDPWR.n132 VDPWR.n16 0.120292
R462 VDPWR.n128 VDPWR.n16 0.120292
R463 VDPWR.n128 VDPWR.n127 0.120292
R464 VDPWR.n127 VDPWR.n19 0.120292
R465 VDPWR.n123 VDPWR.n19 0.120292
R466 VDPWR.n123 VDPWR.n122 0.120292
R467 VDPWR.n122 VDPWR.n121 0.120292
R468 VDPWR.n44 VDPWR.n43 0.120292
R469 VDPWR.n44 VDPWR.n37 0.120292
R470 VDPWR.n37 VDPWR.n36 0.120292
R471 VDPWR.n49 VDPWR.n36 0.120292
R472 VDPWR.n50 VDPWR.n49 0.120292
R473 VDPWR.n51 VDPWR.n50 0.120292
R474 VDPWR.n51 VDPWR.n33 0.120292
R475 VDPWR.n56 VDPWR.n33 0.120292
R476 VDPWR.n57 VDPWR.n56 0.120292
R477 VDPWR.n58 VDPWR.n57 0.120292
R478 VDPWR.n58 VDPWR.n31 0.120292
R479 VDPWR.n31 VDPWR.n29 0.120292
R480 VDPWR.n64 VDPWR.n29 0.120292
R481 VDPWR.n65 VDPWR.n64 0.120292
R482 VDPWR.n66 VDPWR.n65 0.120292
R483 VDPWR.n66 VDPWR.n26 0.120292
R484 VDPWR.n70 VDPWR.n26 0.120292
R485 VDPWR.n111 VDPWR.n72 0.120292
R486 VDPWR.n106 VDPWR.n72 0.120292
R487 VDPWR.n106 VDPWR.n105 0.120292
R488 VDPWR.n105 VDPWR.n104 0.120292
R489 VDPWR.n104 VDPWR.n74 0.120292
R490 VDPWR.n100 VDPWR.n74 0.120292
R491 VDPWR.n100 VDPWR.n99 0.120292
R492 VDPWR.n99 VDPWR.n77 0.120292
R493 VDPWR.n95 VDPWR.n77 0.120292
R494 VDPWR.n95 VDPWR.n94 0.120292
R495 VDPWR.n94 VDPWR.n93 0.120292
R496 VDPWR.n93 VDPWR.n79 0.120292
R497 VDPWR.n88 VDPWR.n79 0.120292
R498 VDPWR.n88 VDPWR.n87 0.120292
R499 VDPWR.n87 VDPWR.n86 0.120292
R500 VDPWR.n354 VDPWR.n353 0.12023
R501 VDPWR.n214 VDPWR.n213 0.12023
R502 VDPWR.n353 VDPWR.n352 0.119565
R503 VDPWR.n213 VDPWR.n212 0.119565
R504 VDPWR.n292 VDPWR.n291 0.118556
R505 VDPWR.n372 VDPWR.n371 0.118451
R506 VDPWR.n269 VDPWR.n268 0.117381
R507 VDPWR.n189 VDPWR.n188 0.117018
R508 VDPWR.n190 VDPWR.n189 0.116571
R509 VDPWR.n352 VDPWR.n351 0.115278
R510 VDPWR.n212 VDPWR.n211 0.115278
R511 VDPWR.n293 VDPWR.n292 0.114758
R512 VDPWR.n255 VDPWR.n254 0.114696
R513 VDPWR.n311 VDPWR.n201 0.114511
R514 VDPWR.n351 VDPWR.n350 0.114352
R515 VDPWR.n211 VDPWR.n210 0.114352
R516 VDPWR.n267 VDPWR.n266 0.114094
R517 VDPWR.n210 VDPWR.n209 0.113756
R518 VDPWR.n350 VDPWR.n349 0.113235
R519 VDPWR.n257 VDPWR.n256 0.113192
R520 VDPWR.n266 VDPWR.n265 0.113154
R521 VDPWR.n256 VDPWR.n255 0.112678
R522 VDPWR.n259 VDPWR.n258 0.112433
R523 VDPWR.n203 VDPWR.n202 0.112207
R524 VDPWR.n191 VDPWR.n190 0.111422
R525 VDPWR.n209 VDPWR.n208 0.111333
R526 VDPWR.n263 VDPWR.n262 0.111285
R527 VDPWR.n348 VDPWR.n347 0.111081
R528 VDPWR.n208 VDPWR.n207 0.111081
R529 VDPWR.n294 VDPWR.n293 0.111077
R530 VDPWR.n349 VDPWR.n348 0.110429
R531 VDPWR.n261 VDPWR.n260 0.110229
R532 VDPWR.n347 VDPWR.n346 0.11011
R533 VDPWR.n258 VDPWR.n257 0.109923
R534 VDPWR.n268 VDPWR.n267 0.10979
R535 VDPWR.n193 VDPWR.n192 0.109555
R536 VDPWR.n337 VDPWR.n336 0.108951
R537 VDPWR.n345 VDPWR.n344 0.108673
R538 VDPWR.n205 VDPWR.n204 0.108673
R539 VDPWR.n207 VDPWR.n206 0.108622
R540 VDPWR.n264 VDPWR.n263 0.108359
R541 VDPWR.n265 VDPWR.n264 0.108286
R542 VDPWR.n260 VDPWR.n259 0.10823
R543 VDPWR.n192 VDPWR.n191 0.107819
R544 VDPWR.n262 VDPWR.n261 0.107643
R545 VDPWR.n346 VDPWR.n345 0.107267
R546 VDPWR.n206 VDPWR.n205 0.107267
R547 VDPWR.n343 VDPWR.n342 0.107106
R548 VDPWR.n295 VDPWR.n294 0.106561
R549 VDPWR.n194 VDPWR.n193 0.105203
R550 VDPWR.n195 VDPWR.n194 0.105131
R551 VDPWR.n338 VDPWR.n337 0.104693
R552 VDPWR.n339 VDPWR.n338 0.104583
R553 VDPWR.n197 VDPWR.n196 0.104583
R554 VDPWR.n196 VDPWR.n195 0.104127
R555 VDPWR.n340 VDPWR.n339 0.103965
R556 VDPWR.n198 VDPWR.n197 0.103965
R557 VDPWR.n341 VDPWR.n340 0.103813
R558 VDPWR.n201 VDPWR.n198 0.103813
R559 VDPWR.n342 VDPWR.n341 0.103788
R560 VDPWR.n344 VDPWR.n343 0.103439
R561 VDPWR.n204 VDPWR.n203 0.103439
R562 VDPWR.n217 VDPWR.n216 0.100519
R563 VDPWR.n147 VDPWR 0.0981562
R564 VDPWR.n43 VDPWR 0.0981562
R565 VDPWR VDPWR.n111 0.0981562
R566 VDPWR.n357 VDPWR.n356 0.0979265
R567 VDPWR.n297 VDPWR.n296 0.0979265
R568 VDPWR.n356 VDPWR.n154 0.0960882
R569 VDPWR.n298 VDPWR.n297 0.0960882
R570 VDPWR.n155 VDPWR.n154 0.0915714
R571 VDPWR.n299 VDPWR.n298 0.0915714
R572 VDPWR.n156 VDPWR.n155 0.088
R573 VDPWR.n300 VDPWR.n299 0.088
R574 VDPWR.n157 VDPWR.n156 0.0855694
R575 VDPWR.n301 VDPWR.n300 0.0855694
R576 VDPWR.n2 VDPWR.n1 0.0849982
R577 VDPWR.n295 VDPWR.n217 0.0844552
R578 VDPWR.n290 VDPWR.n287 0.0832089
R579 VDPWR.n158 VDPWR.n157 0.0820972
R580 VDPWR.n302 VDPWR.n301 0.0820972
R581 VDPWR.n159 VDPWR.n158 0.0792671
R582 VDPWR.n303 VDPWR.n302 0.0792671
R583 VDPWR.n368 VDPWR.n367 0.078657
R584 VDPWR.n304 VDPWR.n303 0.0775548
R585 VDPWR.n160 VDPWR.n159 0.0765135
R586 VDPWR.n253 VDPWR.n2 0.0741301
R587 VDPWR.n161 VDPWR.n160 0.0731351
R588 VDPWR.n253 VDPWR.n252 0.0724178
R589 VDPWR.n305 VDPWR.n304 0.0721667
R590 VDPWR.n162 VDPWR.n161 0.0705
R591 VDPWR.n306 VDPWR.n305 0.0705
R592 VDPWR.n252 VDPWR.n251 0.0688333
R593 VDPWR.n163 VDPWR.n162 0.0679342
R594 VDPWR.n307 VDPWR.n306 0.0679342
R595 VDPWR.n311 VDPWR.n310 0.0676642
R596 VDPWR.n251 VDPWR.n250 0.0655
R597 VDPWR.n164 VDPWR.n163 0.0646447
R598 VDPWR.n308 VDPWR.n307 0.0646447
R599 VDPWR.n250 VDPWR.n249 0.0646447
R600 VDPWR.n165 VDPWR.n164 0.063
R601 VDPWR.n309 VDPWR.n308 0.063
R602 VDPWR.n121 VDPWR 0.0603958
R603 VDPWR.n23 VDPWR 0.0603958
R604 VDPWR.n40 VDPWR 0.0603958
R605 VDPWR.n42 VDPWR 0.0603958
R606 VDPWR VDPWR.n70 0.0603958
R607 VDPWR.n71 VDPWR 0.0603958
R608 VDPWR.n113 VDPWR 0.0603958
R609 VDPWR VDPWR.n112 0.0603958
R610 VDPWR.n249 VDPWR.n248 0.0597105
R611 VDPWR.n166 VDPWR.n165 0.0589416
R612 VDPWR.n310 VDPWR.n309 0.0589416
R613 VDPWR.n248 VDPWR.n247 0.0581923
R614 VDPWR.n167 VDPWR.n166 0.057462
R615 VDPWR.n8 VDPWR 0.0573182
R616 VDPWR.n226 VDPWR 0.0573182
R617 VDPWR.n223 VDPWR 0.0573182
R618 VDPWR.n178 VDPWR 0.0573182
R619 VDPWR.n174 VDPWR 0.0573182
R620 VDPWR.n153 VDPWR 0.0573182
R621 VDPWR.n361 VDPWR 0.0573182
R622 VDPWR.n364 VDPWR 0.0573182
R623 VDPWR.n200 VDPWR 0.0573182
R624 VDPWR.n289 VDPWR 0.0573182
R625 VDPWR.n247 VDPWR.n246 0.0556948
R626 VDPWR.n168 VDPWR.n167 0.0542975
R627 VDPWR.n169 VDPWR.n168 0.0527152
R628 VDPWR.n313 VDPWR.n312 0.0527152
R629 VDPWR.n246 VDPWR.n245 0.0527152
R630 VDPWR.n4 VDPWR 0.0505
R631 VDPWR.n231 VDPWR 0.0505
R632 VDPWR.n279 VDPWR 0.0505
R633 VDPWR.n229 VDPWR 0.0505
R634 VDPWR.n233 VDPWR 0.0505
R635 VDPWR VDPWR.n373 0.0505
R636 VDPWR.n245 VDPWR.n244 0.0495506
R637 VDPWR.n170 VDPWR.n169 0.0483395
R638 VDPWR.n314 VDPWR.n313 0.0483395
R639 VDPWR.n244 VDPWR.n243 0.0479684
R640 VDPWR.n171 VDPWR.n170 0.047375
R641 VDPWR.n315 VDPWR.n314 0.047375
R642 VDPWR.n312 VDPWR.n311 0.0472033
R643 VDPWR.n172 VDPWR.n171 0.0463861
R644 VDPWR.n316 VDPWR.n315 0.0452531
R645 VDPWR.n243 VDPWR.n242 0.0452531
R646 VDPWR.n242 VDPWR.n241 0.0426875
R647 VDPWR.n317 VDPWR.n316 0.0416585
R648 VDPWR.n175 VDPWR.n172 0.0406786
R649 VDPWR.n372 VDPWR.n1 0.039507
R650 VDPWR.n241 VDPWR.n240 0.0390802
R651 VDPWR.n319 VDPWR.n318 0.0386098
R652 VDPWR.n318 VDPWR.n317 0.0386098
R653 VDPWR.n240 VDPWR.n239 0.0386098
R654 VDPWR VDPWR.n23 0.0382604
R655 VDPWR VDPWR.n40 0.0382604
R656 VDPWR VDPWR.n71 0.0382604
R657 VDPWR.n113 VDPWR 0.0382604
R658 VDPWR.n239 VDPWR.n238 0.035561
R659 VDPWR.n320 VDPWR.n319 0.0351386
R660 VDPWR.n275 VDPWR.n274 0.0350681
R661 VDPWR.n238 VDPWR.n237 0.0325122
R662 VDPWR.n321 VDPWR.n320 0.0321265
R663 VDPWR.n237 VDPWR.n236 0.0306205
R664 VDPWR.n322 VDPWR.n321 0.0302619
R665 VDPWR.n236 VDPWR.n235 0.0276084
R666 VDPWR.n323 VDPWR.n322 0.0272857
R667 VDPWR.n324 VDPWR.n323 0.0257976
R668 VDPWR.n274 VDPWR.n235 0.0257976
R669 VDPWR.n333 VDPWR.n332 0.0244583
R670 VDPWR.n325 VDPWR.n324 0.0243095
R671 VDPWR.n334 VDPWR.n333 0.0239375
R672 VDPWR.n335 VDPWR.n175 0.0227865
R673 VDPWR VDPWR.n42 0.0226354
R674 VDPWR.n112 VDPWR 0.0226354
R675 VDPWR.n149 VDPWR 0.0224072
R676 VDPWR.n326 VDPWR.n325 0.0210882
R677 VDPWR.n327 VDPWR.n326 0.0198452
R678 VDPWR.n328 VDPWR.n327 0.0166765
R679 VDPWR.n329 VDPWR.n328 0.0152059
R680 VDPWR.n273 VDPWR.n234 0.0131488
R681 VDPWR.n330 VDPWR.n329 0.0121279
R682 VDPWR.n331 VDPWR.n330 0.0107941
R683 VDPWR.n359 VDPWR.n358 0.0104434
R684 VDPWR.n332 VDPWR.n331 0.00785294
R685 VDPWR.n291 VDPWR.n290 0.00590164
R686 VGND.n336 VGND.n151 171881
R687 VGND.n342 VGND.n341 156443
R688 VGND.n337 VGND.t61 151322
R689 VGND.n164 VGND.n163 130569
R690 VGND.n368 VGND.n367 130542
R691 VGND.n326 VGND.n162 49690.4
R692 VGND.n370 VGND.n369 48636.9
R693 VGND.n333 VGND.n164 45450.3
R694 VGND.n368 VGND.n75 44132.5
R695 VGND.n163 VGND.n64 44106
R696 VGND.n419 VGND.n65 43377.2
R697 VGND.t67 VGND.n64 31560.8
R698 VGND.n111 VGND.n75 30151.8
R699 VGND.n419 VGND.n64 29891.4
R700 VGND.n108 VGND.n75 29891.4
R701 VGND.n327 VGND.t63 18687.3
R702 VGND.n333 VGND.n151 16600.2
R703 VGND.n375 VGND.n68 16072.7
R704 VGND.n159 VGND.n150 14081.5
R705 VGND.n326 VGND.n63 13406.4
R706 VGND.n327 VGND.n325 13301.5
R707 VGND.n74 VGND.n71 12272.6
R708 VGND.n157 VGND.n71 12077.4
R709 VGND.n333 VGND.n161 11373.6
R710 VGND.n163 VGND.n65 10649.3
R711 VGND.n369 VGND.n368 10649.2
R712 VGND.n333 VGND.n162 8289.38
R713 VGND.n69 VGND.t72 6802.38
R714 VGND.n160 VGND.n65 6127.89
R715 VGND.n371 VGND.n71 5980.78
R716 VGND.n327 VGND 5326.64
R717 VGND.n374 VGND.n68 4541.14
R718 VGND.n66 VGND.n63 4245.54
R719 VGND.n375 VGND.n69 4122.66
R720 VGND.n330 VGND.n329 4044.64
R721 VGND.n330 VGND.t0 3942.35
R722 VGND.n372 VGND.n371 3902.89
R723 VGND.n371 VGND.n370 3517.03
R724 VGND.n333 VGND.n332 3472.59
R725 VGND.n341 VGND.n340 3392.44
R726 VGND.n97 VGND.n68 3164.24
R727 VGND.n100 VGND.n69 3164.24
R728 VGND.n159 VGND.n74 2758.39
R729 VGND.n335 VGND.n333 2554.5
R730 VGND.n340 VGND.t21 2448.45
R731 VGND.n327 VGND 2380.9
R732 VGND.n159 VGND.n158 2252.33
R733 VGND.n333 VGND.n160 2096.68
R734 VGND.n420 VGND.n63 1953.47
R735 VGND.n342 VGND.n151 1821.62
R736 VGND.n73 VGND.t35 1524.56
R737 VGND.n419 VGND.n418 1397.72
R738 VGND.n325 VGND.t19 1303.08
R739 VGND.n370 VGND.n72 1261.32
R740 VGND.n156 VGND.n155 1170
R741 VGND.n154 VGND.n153 1170
R742 VGND.n335 VGND.n334 1170
R743 VGND.n339 VGND.n338 1170
R744 VGND.n325 VGND.n324 1170
R745 VGND.n110 VGND.n109 1170
R746 VGND.n113 VGND.n112 1170
R747 VGND.n106 VGND.n72 1170
R748 VGND.n366 VGND.n365 1170
R749 VGND.n344 VGND.n343 1170
R750 VGND.n167 VGND.n166 1170
R751 VGND.n332 VGND.n331 1170
R752 VGND.n421 VGND.n420 1170
R753 VGND.n377 VGND.n376 1170
R754 VGND.n102 VGND.n70 1170
R755 VGND.n374 VGND.n373 1170
R756 VGND.n104 VGND.n73 1170
R757 VGND.n329 VGND.n328 1170
R758 VGND.n366 VGND.t17 1134.17
R759 VGND.n158 VGND.n63 1052.01
R760 VGND.t52 VGND.n342 876.702
R761 VGND.t9 VGND.n164 844.357
R762 VGND.n150 VGND.n76 843.24
R763 VGND.t15 VGND.n111 753.322
R764 VGND.n419 VGND.n66 747.253
R765 VGND.t61 VGND.n154 713.466
R766 VGND.n108 VGND.t37 696.106
R767 VGND.n340 VGND.n156 646.26
R768 VGND.t48 VGND.n419 629.832
R769 VGND.n323 VGND.n168 595.942
R770 VGND.n323 VGND.n322 595.942
R771 VGND.n111 VGND.n110 585.742
R772 VGND.n112 VGND.n108 546.058
R773 VGND.t21 VGND.n339 508.485
R774 VGND.n333 VGND.n330 493.118
R775 VGND.n66 VGND.t13 467.337
R776 VGND.n329 VGND.t67 380.034
R777 VGND.n167 VGND.n161 333.548
R778 VGND.t76 VGND.n375 302.156
R779 VGND.n109 VGND.t18 282.339
R780 VGND.n102 VGND.t57 282.339
R781 VGND.n373 VGND.t71 282.339
R782 VGND.n334 VGND.t80 282.339
R783 VGND.n344 VGND.t53 282.339
R784 VGND.n365 VGND.t45 282.339
R785 VGND.n338 VGND.t22 282.339
R786 VGND.n100 VGND.t55 282.339
R787 VGND.n104 VGND.t36 282.339
R788 VGND.n106 VGND.t38 282.339
R789 VGND.n113 VGND.t16 282.339
R790 VGND.n377 VGND.t77 282.339
R791 VGND.n421 VGND.t49 282.339
R792 VGND.n328 VGND.t68 282.339
R793 VGND.n155 VGND.t51 282.339
R794 VGND.n153 VGND.t62 282.339
R795 VGND.n166 VGND.t8 282.339
R796 VGND.n331 VGND.t10 282.339
R797 VGND.n324 VGND.t20 282.339
R798 VGND.n418 VGND.t14 282.339
R799 VGND.n97 VGND.t73 282.339
R800 VGND.n332 VGND.t9 266.457
R801 VGND.n247 VGND.t27 251
R802 VGND.n214 VGND.t31 251
R803 VGND.n302 VGND.t5 251
R804 VGND.n336 VGND.t79 248.936
R805 VGND.n234 VGND.t75 243.028
R806 VGND.n201 VGND.t43 243.028
R807 VGND.n315 VGND.t47 243.028
R808 VGND.n69 VGND.t54 236.923
R809 VGND.n327 VGND.n63 219.505
R810 VGND.n249 VGND.n174 218.506
R811 VGND.n188 VGND.n187 218.506
R812 VGND.n270 VGND.n269 218.506
R813 VGND.n370 VGND.n73 212.281
R814 VGND.n255 VGND.n171 200.201
R815 VGND.n185 VGND.n184 200.201
R816 VGND.n273 VGND.n272 200.201
R817 VGND.n183 VGND.n182 199.739
R818 VGND.n197 VGND.n196 199.739
R819 VGND.n261 VGND.n260 199.739
R820 VGND.n240 VGND.n178 199.53
R821 VGND.n207 VGND.n192 199.53
R822 VGND.n309 VGND.n265 199.53
R823 VGND.n372 VGND.n70 199.089
R824 VGND.n339 VGND.n337 190.542
R825 VGND.t79 VGND.n335 187.446
R826 VGND.n157 VGND.t56 183.096
R827 VGND.n112 VGND.t15 170.459
R828 VGND.n420 VGND.t48 169.868
R829 VGND.n110 VGND.t17 166.094
R830 VGND.n330 VGND.n327 165.339
R831 VGND.n333 VGND.t7 159.488
R832 VGND.t37 VGND.n72 158.115
R833 VGND.n341 VGND.n154 144.5
R834 VGND.t56 VGND.n70 140.434
R835 VGND.n161 VGND.t50 132.02
R836 VGND.t2 VGND.n162 128.904
R837 VGND.n343 VGND.t52 124.144
R838 VGND.t7 VGND.n167 122.326
R839 VGND.n375 VGND.t70 120.314
R840 VGND.n376 VGND.t76 111.326
R841 VGND.n158 VGND.n157 104.849
R842 VGND VGND.t40 102.412
R843 VGND.t50 VGND.n156 101.258
R844 VGND.n367 VGND.n76 100.996
R845 VGND.t42 VGND.n326 94.8614
R846 VGND.t24 VGND.t58 93.0774
R847 VGND.t70 VGND.n374 92.2804
R848 VGND.t72 VGND.n68 82.4085
R849 VGND.n178 VGND.t81 74.8666
R850 VGND.n192 VGND.t59 74.8666
R851 VGND.n265 VGND.t12 74.8666
R852 VGND.n171 VGND.t26 54.2862
R853 VGND.n184 VGND.t34 54.2862
R854 VGND.n272 VGND.t1 54.2862
R855 VGND.n367 VGND.n366 46.6396
R856 VGND VGND.t65 45.7764
R857 VGND.n369 VGND.n74 45.2738
R858 VGND.n343 VGND.n150 40.8576
R859 VGND.n178 VGND.t78 40.0005
R860 VGND.n192 VGND.t25 40.0005
R861 VGND.n265 VGND.t39 40.0005
R862 VGND.n182 VGND.t23 38.5719
R863 VGND.n182 VGND.t60 38.5719
R864 VGND.n196 VGND.t46 38.5719
R865 VGND.n196 VGND.t64 38.5719
R866 VGND.n260 VGND.t29 38.5719
R867 VGND.n260 VGND.t41 38.5719
R868 VGND.n376 VGND.n63 36.639
R869 VGND.n250 VGND.n172 34.6358
R870 VGND.n254 VGND.n172 34.6358
R871 VGND.n242 VGND.n241 34.6358
R872 VGND.n242 VGND.n176 34.6358
R873 VGND.n246 VGND.n176 34.6358
R874 VGND.n235 VGND.n180 34.6358
R875 VGND.n239 VGND.n180 34.6358
R876 VGND.n219 VGND.n218 34.6358
R877 VGND.n220 VGND.n219 34.6358
R878 VGND.n209 VGND.n208 34.6358
R879 VGND.n209 VGND.n190 34.6358
R880 VGND.n213 VGND.n190 34.6358
R881 VGND.n202 VGND.n194 34.6358
R882 VGND.n206 VGND.n194 34.6358
R883 VGND.n314 VGND.n263 34.6358
R884 VGND.n310 VGND.n263 34.6358
R885 VGND.n308 VGND.n266 34.6358
R886 VGND.n304 VGND.n266 34.6358
R887 VGND.n304 VGND.n303 34.6358
R888 VGND.n298 VGND.n297 34.6358
R889 VGND.n297 VGND.n296 34.6358
R890 VGND.n249 VGND.n248 32.7534
R891 VGND.n215 VGND.n188 32.7534
R892 VGND.n301 VGND.n270 32.7534
R893 VGND.n248 VGND.n247 31.2476
R894 VGND.n215 VGND.n214 31.2476
R895 VGND.n302 VGND.n301 31.2476
R896 VGND.n240 VGND.n239 30.8711
R897 VGND.n207 VGND.n206 30.8711
R898 VGND.n310 VGND.n309 30.8711
R899 VGND.n235 VGND.n234 27.4829
R900 VGND.n202 VGND.n201 27.4829
R901 VGND.n315 VGND.n314 27.4829
R902 VGND.t4 VGND.t11 27.1458
R903 VGND.n171 VGND.t30 25.9346
R904 VGND.n184 VGND.t6 25.9346
R905 VGND.n272 VGND.t74 25.9346
R906 VGND.n375 VGND.n372 25.8467
R907 VGND.t63 VGND.t24 25.3851
R908 VGND.n174 VGND.t82 24.9236
R909 VGND.n174 VGND.t28 24.9236
R910 VGND.n187 VGND.t66 24.9236
R911 VGND.n187 VGND.t33 24.9236
R912 VGND.n269 VGND.t69 24.9236
R913 VGND.n269 VGND.t3 24.9236
R914 VGND.n256 VGND.n169 23.7181
R915 VGND.n255 VGND.n254 23.7181
R916 VGND.n229 VGND.n228 23.7181
R917 VGND.n225 VGND.n224 23.7181
R918 VGND.n220 VGND.n185 23.7181
R919 VGND.n321 VGND.n320 23.7181
R920 VGND.n296 VGND.n273 23.7181
R921 VGND.n233 VGND.n183 22.9652
R922 VGND.n234 VGND.n233 22.9652
R923 VGND.n200 VGND.n197 22.9652
R924 VGND.n201 VGND.n200 22.9652
R925 VGND.n316 VGND.n261 22.9652
R926 VGND.n316 VGND.n315 22.9652
R927 VGND.n247 VGND.n246 22.2123
R928 VGND.n214 VGND.n213 22.2123
R929 VGND.n303 VGND.n302 22.2123
R930 VGND.n256 VGND.n255 21.4593
R931 VGND.n229 VGND.n183 21.4593
R932 VGND.n224 VGND.n185 21.4593
R933 VGND.n320 VGND.n261 21.4593
R934 VGND.n105 VGND.n103 20.9274
R935 VGND.t2 VGND.t0 19.8983
R936 VGND.t2 VGND.n323 19.7425
R937 VGND.n346 VGND.n149 17.0502
R938 VGND.n160 VGND.n159 14.7835
R939 VGND.n378 VGND.n377 13.3141
R940 VGND.n422 VGND.n421 13.3141
R941 VGND.n328 VGND.n40 13.3141
R942 VGND.n155 VGND.n2 13.3141
R943 VGND.n153 VGND.n152 13.3141
R944 VGND.n166 VGND.n165 13.3141
R945 VGND.n331 VGND.n20 13.3141
R946 VGND.n324 VGND.n42 13.3141
R947 VGND.n418 VGND.n417 13.3141
R948 VGND.n98 VGND.n97 13.3141
R949 VGND VGND.n102 13.2586
R950 VGND.n373 VGND 13.2586
R951 VGND VGND.n344 13.2586
R952 VGND.n365 VGND 13.2586
R953 VGND.n334 VGND 13.2586
R954 VGND.n338 VGND 13.2586
R955 VGND VGND.n100 13.2586
R956 VGND VGND.n104 13.2586
R957 VGND VGND.n106 13.2586
R958 VGND VGND.n113 13.2586
R959 VGND.n109 VGND 13.2586
R960 VGND VGND.n293 11.784
R961 VGND VGND.n149 10.8878
R962 VGND.n241 VGND.n240 10.5417
R963 VGND.n208 VGND.n207 10.5417
R964 VGND.n309 VGND.n308 10.5417
R965 VGND.n487 VGND.n486 9.52816
R966 VGND.n488 VGND 9.46719
R967 VGND.n296 VGND.n295 9.3005
R968 VGND.n297 VGND.n271 9.3005
R969 VGND.n299 VGND.n298 9.3005
R970 VGND.n301 VGND.n300 9.3005
R971 VGND.n302 VGND.n268 9.3005
R972 VGND.n303 VGND.n267 9.3005
R973 VGND.n305 VGND.n304 9.3005
R974 VGND.n306 VGND.n266 9.3005
R975 VGND.n308 VGND.n307 9.3005
R976 VGND.n309 VGND.n264 9.3005
R977 VGND.n311 VGND.n310 9.3005
R978 VGND.n312 VGND.n263 9.3005
R979 VGND.n314 VGND.n313 9.3005
R980 VGND.n315 VGND.n262 9.3005
R981 VGND.n317 VGND.n316 9.3005
R982 VGND.n318 VGND.n261 9.3005
R983 VGND.n320 VGND.n319 9.3005
R984 VGND.n321 VGND.n259 9.3005
R985 VGND.n200 VGND.n199 9.3005
R986 VGND.n201 VGND.n195 9.3005
R987 VGND.n203 VGND.n202 9.3005
R988 VGND.n204 VGND.n194 9.3005
R989 VGND.n206 VGND.n205 9.3005
R990 VGND.n207 VGND.n193 9.3005
R991 VGND.n208 VGND.n191 9.3005
R992 VGND.n210 VGND.n209 9.3005
R993 VGND.n211 VGND.n190 9.3005
R994 VGND.n213 VGND.n212 9.3005
R995 VGND.n214 VGND.n189 9.3005
R996 VGND.n216 VGND.n215 9.3005
R997 VGND.n218 VGND.n217 9.3005
R998 VGND.n219 VGND.n186 9.3005
R999 VGND.n221 VGND.n220 9.3005
R1000 VGND.n222 VGND.n185 9.3005
R1001 VGND.n224 VGND.n223 9.3005
R1002 VGND.n226 VGND.n225 9.3005
R1003 VGND.n228 VGND.n227 9.3005
R1004 VGND.n230 VGND.n229 9.3005
R1005 VGND.n231 VGND.n183 9.3005
R1006 VGND.n233 VGND.n232 9.3005
R1007 VGND.n234 VGND.n181 9.3005
R1008 VGND.n236 VGND.n235 9.3005
R1009 VGND.n237 VGND.n180 9.3005
R1010 VGND.n239 VGND.n238 9.3005
R1011 VGND.n240 VGND.n179 9.3005
R1012 VGND.n241 VGND.n177 9.3005
R1013 VGND.n243 VGND.n242 9.3005
R1014 VGND.n244 VGND.n176 9.3005
R1015 VGND.n246 VGND.n245 9.3005
R1016 VGND.n247 VGND.n175 9.3005
R1017 VGND.n248 VGND.n173 9.3005
R1018 VGND.n251 VGND.n250 9.3005
R1019 VGND.n252 VGND.n172 9.3005
R1020 VGND.n254 VGND.n253 9.3005
R1021 VGND.n255 VGND.n170 9.3005
R1022 VGND.n257 VGND.n256 9.3005
R1023 VGND.n258 VGND.n169 9.3005
R1024 VGND.n99 VGND.n98 9.16992
R1025 VGND.n103 VGND 8.69654
R1026 VGND.n379 VGND.n378 8.60727
R1027 VGND.n345 VGND 8.50779
R1028 VGND.n380 VGND.n379 8.47715
R1029 VGND.n152 VGND.n1 7.73586
R1030 VGND.n101 VGND 7.66873
R1031 VGND.t40 VGND.t4 7.40375
R1032 VGND VGND.n364 7.24133
R1033 VGND.n417 VGND.n416 7.18609
R1034 VGND.n198 VGND.n197 7.12576
R1035 VGND.n294 VGND.n273 7.12063
R1036 VGND.n487 VGND.n2 6.8256
R1037 VGND VGND.n67 6.67637
R1038 VGND.n165 VGND.n3 6.61112
R1039 VGND.n423 VGND.n422 6.60276
R1040 VGND VGND.n96 6.5915
R1041 VGND.n114 VGND 6.55995
R1042 VGND.n225 VGND.n168 6.367
R1043 VGND.n322 VGND.n321 6.367
R1044 VGND.n322 VGND.n169 6.367
R1045 VGND.n228 VGND.n168 6.367
R1046 VGND.n105 VGND 6.30778
R1047 VGND.n467 VGND.n20 6.21471
R1048 VGND.n107 VGND 6.20286
R1049 VGND.n444 VGND.n42 6.13644
R1050 VGND.n447 VGND.n40 5.99894
R1051 VGND.n282 VGND.n0 4.70536
R1052 VGND.t58 VGND.t32 4.23127
R1053 VGND.n379 VGND.n67 3.52675
R1054 VGND.n0 VGND 3.44325
R1055 VGND.n491 VGND 3.36335
R1056 VGND.t65 VGND.t42 3.3096
R1057 VGND.n107 VGND.n105 2.92676
R1058 VGND.n488 VGND.n487 2.38171
R1059 VGND VGND.n491 2.34667
R1060 VGND.n337 VGND.n336 2.10058
R1061 VGND.n76 VGND.t44 1.91332
R1062 VGND.n250 VGND.n249 1.88285
R1063 VGND.n218 VGND.n188 1.88285
R1064 VGND.n298 VGND.n270 1.88285
R1065 VGND.n103 VGND.n101 1.59945
R1066 VGND.n114 VGND.n107 1.28972
R1067 VGND.t11 VGND.t2 1.23438
R1068 VGND.n101 VGND.n99 1.05629
R1069 VGND.n489 VGND.n488 0.952529
R1070 VGND.n99 VGND.n67 0.951875
R1071 VGND.n149 VGND.n1 0.752727
R1072 VGND.n115 VGND.n114 0.663554
R1073 VGND.n490 VGND.n489 0.544604
R1074 VGND.n446 VGND.n445 0.457033
R1075 VGND.n274 uo_out[4] 0.39812
R1076 VGND.n444 VGND.n443 0.297375
R1077 VGND.n274 uo_out[5] 0.2684
R1078 VGND.n275 uo_out[6] 0.2684
R1079 VGND.n276 uo_out[7] 0.2684
R1080 VGND.n277 uio_out[0] 0.2684
R1081 VGND.n278 uio_out[1] 0.2684
R1082 VGND.n279 uio_out[2] 0.2684
R1083 VGND.n280 uio_out[3] 0.2684
R1084 VGND.n281 uio_out[4] 0.2684
R1085 VGND.n292 uio_out[5] 0.2684
R1086 VGND.n291 uio_out[6] 0.2684
R1087 VGND.n290 uio_out[7] 0.2684
R1088 VGND.n289 uio_oe[0] 0.2684
R1089 VGND.n288 uio_oe[1] 0.2684
R1090 VGND.n287 uio_oe[2] 0.2684
R1091 VGND.n286 uio_oe[3] 0.2684
R1092 VGND.n285 uio_oe[4] 0.2684
R1093 VGND.n284 uio_oe[5] 0.2684
R1094 VGND.n283 uio_oe[6] 0.2684
R1095 VGND.n282 uio_oe[7] 0.2684
R1096 VGND.n443 VGND.n442 0.240747
R1097 VGND.n132 VGND.n79 0.232444
R1098 VGND.n442 VGND.n441 0.201889
R1099 VGND.n441 VGND.n440 0.183192
R1100 VGND.n486 VGND.n485 0.181207
R1101 VGND.n116 VGND.n115 0.177735
R1102 VGND.n416 VGND.n380 0.15732
R1103 VGND.n347 VGND.n346 0.155253
R1104 VGND.n294 VGND 0.152603
R1105 VGND.n133 VGND.n132 0.152388
R1106 VGND.n295 VGND.n294 0.148519
R1107 VGND.n439 VGND.n438 0.145639
R1108 VGND.n468 VGND.n467 0.14536
R1109 VGND.n440 VGND.n439 0.14425
R1110 VGND.n199 VGND.n198 0.143396
R1111 VGND.n442 VGND.n43 0.135917
R1112 VGND.n443 VGND.n41 0.135115
R1113 VGND.n440 VGND.n45 0.134528
R1114 VGND.n441 VGND.n44 0.133742
R1115 VGND.n445 VGND.n444 0.133539
R1116 VGND.n439 VGND.n46 0.133139
R1117 VGND.n438 VGND.n47 0.133139
R1118 VGND.n437 VGND.n48 0.13175
R1119 VGND.n117 VGND.n94 0.131182
R1120 VGND.n434 VGND.n51 0.131118
R1121 VGND.n436 VGND.n49 0.131056
R1122 VGND.n435 VGND.n50 0.130361
R1123 VGND.n275 VGND.n274 0.13022
R1124 VGND.n276 VGND.n275 0.13022
R1125 VGND.n277 VGND.n276 0.13022
R1126 VGND.n278 VGND.n277 0.13022
R1127 VGND.n279 VGND.n278 0.13022
R1128 VGND.n280 VGND.n279 0.13022
R1129 VGND.n281 VGND.n280 0.13022
R1130 VGND.n292 VGND.n291 0.13022
R1131 VGND.n291 VGND.n290 0.13022
R1132 VGND.n290 VGND.n289 0.13022
R1133 VGND.n289 VGND.n288 0.13022
R1134 VGND.n288 VGND.n287 0.13022
R1135 VGND.n287 VGND.n286 0.13022
R1136 VGND.n286 VGND.n285 0.13022
R1137 VGND.n285 VGND.n284 0.13022
R1138 VGND.n284 VGND.n283 0.13022
R1139 VGND.n283 VGND.n282 0.13022
R1140 VGND.n119 VGND.n92 0.129761
R1141 VGND.n430 VGND.n55 0.129761
R1142 VGND.n116 VGND.n95 0.129713
R1143 VGND.n433 VGND.n52 0.129713
R1144 VGND.n120 VGND.n91 0.128341
R1145 VGND.n118 VGND.n93 0.128309
R1146 VGND.n431 VGND.n54 0.128309
R1147 VGND.n432 VGND.n53 0.128278
R1148 VGND.n125 VGND.n86 0.12768
R1149 VGND.n123 VGND.n88 0.127655
R1150 VGND.n121 VGND.n90 0.127631
R1151 VGND.n448 VGND.n39 0.127631
R1152 VGND.n428 VGND.n57 0.127631
R1153 VGND.n126 VGND.n85 0.126953
R1154 VGND.n124 VGND.n87 0.126937
R1155 VGND.n122 VGND.n89 0.12692
R1156 VGND.n449 VGND.n38 0.12692
R1157 VGND.n427 VGND.n58 0.12692
R1158 VGND.n429 VGND.n56 0.126904
R1159 VGND.n481 VGND.n6 0.126368
R1160 VGND.n347 VGND.n148 0.126345
R1161 VGND.n349 VGND.n146 0.126333
R1162 VGND.n351 VGND.n144 0.126322
R1163 VGND.n353 VGND.n142 0.126312
R1164 VGND.n131 VGND.n80 0.126244
R1165 VGND.n452 VGND.n35 0.126218
R1166 VGND.n424 VGND.n61 0.126218
R1167 VGND.n450 VGND.n37 0.12621
R1168 VGND.n426 VGND.n59 0.12621
R1169 VGND.n127 VGND.n84 0.1255
R1170 VGND.n128 VGND.n83 0.1255
R1171 VGND.n129 VGND.n82 0.1255
R1172 VGND.n358 VGND.n137 0.1255
R1173 VGND.n356 VGND.n139 0.1255
R1174 VGND.n348 VGND.n147 0.1255
R1175 VGND.n455 VGND.n32 0.1255
R1176 VGND.n454 VGND.n33 0.1255
R1177 VGND.n453 VGND.n34 0.1255
R1178 VGND.n451 VGND.n36 0.1255
R1179 VGND.n425 VGND.n60 0.1255
R1180 VGND.n389 VGND.n62 0.1255
R1181 VGND.n391 VGND.n390 0.1255
R1182 VGND.n392 VGND.n388 0.1255
R1183 VGND.n130 VGND.n81 0.124765
R1184 VGND.n458 VGND.n29 0.124765
R1185 VGND.n397 VGND.n396 0.124765
R1186 VGND.n364 VGND.n363 0.124747
R1187 VGND.n361 VGND.n134 0.124738
R1188 VGND.n359 VGND.n136 0.124728
R1189 VGND.n355 VGND.n140 0.124709
R1190 VGND.n473 VGND.n14 0.124688
R1191 VGND.n475 VGND.n12 0.124678
R1192 VGND.n477 VGND.n10 0.124667
R1193 VGND.n480 VGND.n7 0.124655
R1194 VGND.n479 VGND.n8 0.124655
R1195 VGND.n482 VGND.n5 0.124644
R1196 VGND.n456 VGND.n31 0.124047
R1197 VGND.n394 VGND.n393 0.124047
R1198 VGND.n460 VGND.n27 0.124012
R1199 VGND.n400 VGND.n399 0.124012
R1200 VGND.n362 VGND.n78 0.123994
R1201 VGND.n462 VGND.n25 0.123994
R1202 VGND.n403 VGND.n402 0.123994
R1203 VGND.n360 VGND.n135 0.123976
R1204 VGND.n412 VGND.n411 0.123938
R1205 VGND.n354 VGND.n141 0.123918
R1206 VGND.n470 VGND.n17 0.123918
R1207 VGND.n415 VGND.n414 0.123918
R1208 VGND.n352 VGND.n143 0.123897
R1209 VGND.n350 VGND.n145 0.123877
R1210 VGND.n478 VGND.n9 0.123833
R1211 VGND.n469 VGND.n468 0.123779
R1212 VGND.n457 VGND.n30 0.12332
R1213 VGND.n395 VGND.n387 0.12332
R1214 VGND.n459 VGND.n28 0.123294
R1215 VGND.n398 VGND.n386 0.123294
R1216 VGND.n461 VGND.n26 0.123268
R1217 VGND.n401 VGND.n385 0.123268
R1218 VGND.n463 VGND.n24 0.123241
R1219 VGND.n404 VGND.n384 0.123241
R1220 VGND.n407 VGND.n383 0.123213
R1221 VGND.n357 VGND.n138 0.123185
R1222 VGND.n410 VGND.n382 0.123185
R1223 VGND.n471 VGND.n16 0.123127
R1224 VGND.n464 VGND.n23 0.122488
R1225 VGND.n406 VGND.n405 0.122488
R1226 VGND.n409 VGND.n408 0.122451
R1227 VGND.n472 VGND.n15 0.122335
R1228 VGND.n474 VGND.n13 0.122295
R1229 VGND.n476 VGND.n11 0.122253
R1230 VGND.n469 VGND.n18 0.121642
R1231 VGND.n413 VGND.n381 0.121642
R1232 VGND.n293 VGND.n292 0.12129
R1233 VGND.n438 VGND.n437 0.120386
R1234 VGND.n199 VGND.n195 0.120292
R1235 VGND.n203 VGND.n195 0.120292
R1236 VGND.n204 VGND.n203 0.120292
R1237 VGND.n205 VGND.n204 0.120292
R1238 VGND.n205 VGND.n193 0.120292
R1239 VGND.n193 VGND.n191 0.120292
R1240 VGND.n210 VGND.n191 0.120292
R1241 VGND.n211 VGND.n210 0.120292
R1242 VGND.n212 VGND.n211 0.120292
R1243 VGND.n212 VGND.n189 0.120292
R1244 VGND.n216 VGND.n189 0.120292
R1245 VGND.n217 VGND.n216 0.120292
R1246 VGND.n217 VGND.n186 0.120292
R1247 VGND.n221 VGND.n186 0.120292
R1248 VGND.n222 VGND.n221 0.120292
R1249 VGND.n223 VGND.n222 0.120292
R1250 VGND.n232 VGND.n231 0.120292
R1251 VGND.n232 VGND.n181 0.120292
R1252 VGND.n236 VGND.n181 0.120292
R1253 VGND.n237 VGND.n236 0.120292
R1254 VGND.n238 VGND.n237 0.120292
R1255 VGND.n238 VGND.n179 0.120292
R1256 VGND.n179 VGND.n177 0.120292
R1257 VGND.n243 VGND.n177 0.120292
R1258 VGND.n244 VGND.n243 0.120292
R1259 VGND.n245 VGND.n244 0.120292
R1260 VGND.n245 VGND.n175 0.120292
R1261 VGND.n175 VGND.n173 0.120292
R1262 VGND.n251 VGND.n173 0.120292
R1263 VGND.n252 VGND.n251 0.120292
R1264 VGND.n253 VGND.n252 0.120292
R1265 VGND.n253 VGND.n170 0.120292
R1266 VGND.n257 VGND.n170 0.120292
R1267 VGND.n318 VGND.n317 0.120292
R1268 VGND.n317 VGND.n262 0.120292
R1269 VGND.n313 VGND.n262 0.120292
R1270 VGND.n313 VGND.n312 0.120292
R1271 VGND.n312 VGND.n311 0.120292
R1272 VGND.n311 VGND.n264 0.120292
R1273 VGND.n307 VGND.n264 0.120292
R1274 VGND.n307 VGND.n306 0.120292
R1275 VGND.n306 VGND.n305 0.120292
R1276 VGND.n305 VGND.n267 0.120292
R1277 VGND.n268 VGND.n267 0.120292
R1278 VGND.n300 VGND.n268 0.120292
R1279 VGND.n300 VGND.n299 0.120292
R1280 VGND.n299 VGND.n271 0.120292
R1281 VGND.n295 VGND.n271 0.120292
R1282 VGND.n484 VGND.n483 0.115369
R1283 VGND.n437 VGND.n436 0.112306
R1284 VGND.n482 VGND.n481 0.111879
R1285 VGND.n483 VGND.n482 0.111186
R1286 VGND.n436 VGND.n435 0.109795
R1287 VGND.n480 VGND.n479 0.108943
R1288 VGND.n132 VGND.n131 0.108833
R1289 VGND.n481 VGND.n480 0.107764
R1290 VGND.n435 VGND.n434 0.107742
R1291 VGND.n479 VGND.n478 0.107535
R1292 VGND.n414 VGND.n380 0.107341
R1293 VGND.n478 VGND.n477 0.106725
R1294 VGND.n348 VGND.n347 0.106074
R1295 VGND.n349 VGND.n348 0.105969
R1296 VGND.n476 VGND.n475 0.1059
R1297 VGND.n350 VGND.n349 0.105163
R1298 VGND.n477 VGND.n476 0.104834
R1299 VGND.n475 VGND.n474 0.104121
R1300 VGND.n474 VGND.n473 0.103867
R1301 VGND.n351 VGND.n350 0.10332
R1302 VGND.n352 VGND.n351 0.10304
R1303 VGND.n118 VGND.n117 0.102984
R1304 VGND.n354 VGND.n353 0.102502
R1305 VGND.n471 VGND.n470 0.102274
R1306 VGND.n473 VGND.n472 0.10217
R1307 VGND.n472 VGND.n471 0.101442
R1308 VGND.n353 VGND.n352 0.101279
R1309 VGND.n411 VGND.n381 0.1005
R1310 VGND.n356 VGND.n355 0.100144
R1311 VGND.n411 VGND.n410 0.0994435
R1312 VGND.n357 VGND.n356 0.099433
R1313 VGND.n355 VGND.n354 0.0992982
R1314 VGND.n470 VGND.n469 0.0991552
R1315 VGND.n415 VGND.n381 0.0991552
R1316 VGND.n21 VGND.n19 0.0981562
R1317 VGND.n231 VGND 0.0981562
R1318 VGND VGND.n318 0.0981562
R1319 VGND.n466 VGND.n465 0.0977932
R1320 VGND.n409 VGND.n383 0.0977932
R1321 VGND.n359 VGND.n358 0.0976284
R1322 VGND.n465 VGND.n464 0.0968228
R1323 VGND.n405 VGND.n383 0.0968228
R1324 VGND.n410 VGND.n409 0.0966929
R1325 VGND.n360 VGND.n359 0.0965648
R1326 VGND.n358 VGND.n357 0.0962384
R1327 VGND.n464 VGND.n463 0.0962186
R1328 VGND.n405 VGND.n404 0.0962186
R1329 VGND.n7 VGND.n6 0.0959861
R1330 VGND.n463 VGND.n462 0.0956231
R1331 VGND.n404 VGND.n403 0.0956231
R1332 VGND.n361 VGND.n360 0.0955348
R1333 VGND.n362 VGND.n361 0.0948777
R1334 VGND.n6 VGND.n5 0.0946781
R1335 VGND.n120 VGND.n119 0.0945657
R1336 VGND.n117 VGND.n116 0.0938949
R1337 VGND.n433 VGND.n432 0.0937672
R1338 VGND.n119 VGND.n118 0.0931452
R1339 VGND.n431 VGND.n430 0.0930016
R1340 VGND.n465 VGND.n22 0.0927256
R1341 VGND.n462 VGND.n461 0.0927181
R1342 VGND.n403 VGND.n385 0.0927181
R1343 VGND.n434 VGND.n433 0.0923627
R1344 VGND.n79 VGND.n77 0.0921667
R1345 VGND.n461 VGND.n460 0.0920855
R1346 VGND.n399 VGND.n385 0.0920855
R1347 VGND.n363 VGND.n362 0.0919467
R1348 VGND.n432 VGND.n431 0.0914722
R1349 VGND.n363 VGND.n133 0.0912494
R1350 VGND.n460 VGND.n459 0.091171
R1351 VGND.n399 VGND.n398 0.091171
R1352 VGND.n121 VGND.n120 0.0904148
R1353 VGND.n8 VGND.n7 0.090027
R1354 VGND.n9 VGND.n8 0.090027
R1355 VGND.n459 VGND.n458 0.0898264
R1356 VGND.n398 VGND.n397 0.0898264
R1357 VGND.n457 VGND.n456 0.0891127
R1358 VGND.n393 VGND.n387 0.0891127
R1359 VGND.n127 VGND.n126 0.0881565
R1360 VGND.n131 VGND.n130 0.0881488
R1361 VGND.n130 VGND.n129 0.0879493
R1362 VGND.n456 VGND.n455 0.0878131
R1363 VGND.n393 VGND.n392 0.0878131
R1364 VGND.n458 VGND.n457 0.0876124
R1365 VGND.n397 VGND.n387 0.0876124
R1366 VGND.n122 VGND.n121 0.0875536
R1367 VGND.n10 VGND.n9 0.0871667
R1368 VGND.n126 VGND.n125 0.0868953
R1369 VGND.n345 VGND.n148 0.0866486
R1370 VGND.n125 VGND.n124 0.0863769
R1371 VGND.n429 VGND.n428 0.0859735
R1372 VGND.n124 VGND.n123 0.0856762
R1373 VGND.n133 VGND.n77 0.085541
R1374 VGND.n11 VGND.n10 0.0855
R1375 VGND.n123 VGND.n122 0.0852048
R1376 VGND.n430 VGND.n429 0.0851591
R1377 VGND.n129 VGND.n128 0.0850588
R1378 VGND.n148 VGND.n147 0.0838333
R1379 VGND.n449 VGND.n448 0.0835966
R1380 VGND.n428 VGND.n427 0.0835966
R1381 VGND.n453 VGND.n452 0.0833636
R1382 VGND.n128 VGND.n127 0.0833488
R1383 VGND.n455 VGND.n454 0.0833488
R1384 VGND.n392 VGND.n391 0.0833488
R1385 VGND.n452 VGND.n451 0.0825455
R1386 VGND.n147 VGND.n146 0.0821667
R1387 VGND.n423 VGND.n62 0.081981
R1388 VGND.n451 VGND.n450 0.0819394
R1389 VGND.n426 VGND.n425 0.0819394
R1390 VGND.n454 VGND.n453 0.0816782
R1391 VGND.n391 VGND.n62 0.0816782
R1392 VGND.n12 VGND.n11 0.0816688
R1393 VGND.n450 VGND.n449 0.0813424
R1394 VGND.n427 VGND.n426 0.0813424
R1395 VGND.n13 VGND.n12 0.0810921
R1396 VGND.n468 VGND.n19 0.0797137
R1397 VGND.n484 VGND.n3 0.0796453
R1398 VGND.n5 VGND.n4 0.0796157
R1399 VGND.n146 VGND.n145 0.0784221
R1400 VGND.n145 VGND.n144 0.0778026
R1401 VGND.n14 VGND.n13 0.0774231
R1402 VGND.n15 VGND.n14 0.0767987
R1403 VGND.n483 VGND.n4 0.0762042
R1404 VGND.n198 VGND 0.0758148
R1405 VGND.n144 VGND.n143 0.074218
R1406 VGND.n143 VGND.n142 0.073552
R1407 VGND.n16 VGND.n15 0.0732848
R1408 VGND.n447 VGND.n446 0.0732142
R1409 VGND.n448 VGND.n447 0.0719286
R1410 VGND.n17 VGND.n16 0.0717025
R1411 VGND.n142 VGND.n141 0.0701203
R1412 VGND.n18 VGND.n17 0.0701203
R1413 VGND.n414 VGND.n413 0.0701203
R1414 VGND.n141 VGND.n140 0.068538
R1415 VGND.n140 VGND.n139 0.0669557
R1416 VGND.n19 VGND.n18 0.066858
R1417 VGND.n413 VGND.n412 0.066858
R1418 VGND.n23 VGND.n22 0.0667809
R1419 VGND.n412 VGND.n382 0.066125
R1420 VGND.n139 VGND.n138 0.0637716
R1421 VGND.n408 VGND.n382 0.0637716
R1422 VGND.n138 VGND.n137 0.063
R1423 VGND.n408 VGND.n407 0.0614756
R1424 VGND.n425 VGND.n424 0.0609482
R1425 VGND.n137 VGND.n136 0.0606852
R1426 VGND.n223 VGND 0.0603958
R1427 VGND.n226 VGND 0.0603958
R1428 VGND.n227 VGND 0.0603958
R1429 VGND.n230 VGND 0.0603958
R1430 VGND VGND.n257 0.0603958
R1431 VGND.n258 VGND 0.0603958
R1432 VGND.n259 VGND 0.0603958
R1433 VGND.n319 VGND 0.0603958
R1434 VGND.n407 VGND.n406 0.0599512
R1435 VGND.n136 VGND.n135 0.0584268
R1436 VGND.n24 VGND.n23 0.0577289
R1437 VGND.n406 VGND.n384 0.0577289
R1438 VGND.n135 VGND.n134 0.0569024
R1439 VGND.n25 VGND.n24 0.0562229
R1440 VGND.n402 VGND.n384 0.0562229
R1441 VGND.n378 VGND 0.0560556
R1442 VGND.n422 VGND 0.0560556
R1443 VGND.n40 VGND 0.0560556
R1444 VGND.n2 VGND 0.0560556
R1445 VGND.n152 VGND 0.0560556
R1446 VGND.n165 VGND 0.0560556
R1447 VGND.n20 VGND 0.0560556
R1448 VGND.n42 VGND 0.0560556
R1449 VGND.n417 VGND 0.0560556
R1450 VGND.n98 VGND 0.0560556
R1451 VGND.n486 VGND.n3 0.0554302
R1452 VGND.n134 VGND.n78 0.0547169
R1453 VGND.n26 VGND.n25 0.0547169
R1454 VGND.n402 VGND.n401 0.0547169
R1455 VGND.n364 VGND.n78 0.0532108
R1456 VGND.n27 VGND.n26 0.0525833
R1457 VGND.n401 VGND.n400 0.0525833
R1458 VGND.n485 VGND.n4 0.0514752
R1459 VGND.n28 VGND.n27 0.0510952
R1460 VGND.n400 VGND.n386 0.0510952
R1461 VGND.n29 VGND.n28 0.0490294
R1462 VGND.n396 VGND.n386 0.0490294
R1463 VGND.n446 VGND.n39 0.0488306
R1464 VGND.n80 VGND.n79 0.046631
R1465 VGND.n466 VGND.n21 0.0461288
R1466 VGND.n81 VGND.n80 0.0460882
R1467 VGND.n30 VGND.n29 0.0460882
R1468 VGND.n396 VGND.n395 0.0460882
R1469 VGND.n31 VGND.n30 0.0455581
R1470 VGND.n395 VGND.n394 0.0455581
R1471 VGND.n82 VGND.n81 0.0446176
R1472 VGND.n32 VGND.n31 0.0441047
R1473 VGND.n394 VGND.n388 0.0441047
R1474 VGND.n84 VGND.n83 0.0411977
R1475 VGND.n83 VGND.n82 0.0411977
R1476 VGND.n33 VGND.n32 0.0411977
R1477 VGND.n34 VGND.n33 0.0411977
R1478 VGND.n390 VGND.n389 0.0411977
R1479 VGND.n390 VGND.n388 0.0411977
R1480 VGND.n346 VGND.n345 0.0401474
R1481 VGND.n85 VGND.n84 0.0382907
R1482 VGND.n485 VGND.n484 0.0381773
R1483 VGND.n35 VGND.n34 0.0378563
R1484 VGND.n389 VGND.n61 0.0378563
R1485 VGND.n86 VGND.n85 0.0368372
R1486 VGND.n36 VGND.n35 0.0364195
R1487 VGND.n61 VGND.n60 0.0364195
R1488 VGND.n364 VGND.n77 0.0353361
R1489 VGND.n416 VGND.n415 0.0353101
R1490 VGND.n87 VGND.n86 0.0349828
R1491 VGND.n37 VGND.n36 0.0345909
R1492 VGND.n60 VGND.n59 0.0345909
R1493 VGND VGND.n226 0.0343542
R1494 VGND.n227 VGND 0.0343542
R1495 VGND VGND.n258 0.0343542
R1496 VGND VGND.n259 0.0343542
R1497 VGND.n88 VGND.n87 0.033546
R1498 VGND.n38 VGND.n37 0.0331705
R1499 VGND.n59 VGND.n58 0.0331705
R1500 VGND.n89 VGND.n88 0.03175
R1501 VGND.n39 VGND.n38 0.03175
R1502 VGND.n58 VGND.n57 0.03175
R1503 VGND.n22 VGND.n21 0.0315583
R1504 VGND.n90 VGND.n89 0.0303295
R1505 VGND.n57 VGND.n56 0.0303295
R1506 VGND.n91 VGND.n90 0.0289091
R1507 VGND.n56 VGND.n55 0.0285899
R1508 VGND.n490 VGND.n0 0.0283721
R1509 VGND.n491 VGND.n490 0.0283721
R1510 VGND.n92 VGND.n91 0.0260682
R1511 VGND.n55 VGND.n54 0.0260682
R1512 VGND.n93 VGND.n92 0.0257809
R1513 VGND.n54 VGND.n53 0.0257809
R1514 VGND.n94 VGND.n93 0.0232273
R1515 VGND.n95 VGND.n94 0.0229719
R1516 VGND.n52 VGND.n51 0.0229719
R1517 VGND.n53 VGND.n52 0.0227222
R1518 VGND VGND.n230 0.0226354
R1519 VGND.n319 VGND 0.0226354
R1520 VGND.n51 VGND.n50 0.0201629
R1521 VGND.n96 VGND.n95 0.0199444
R1522 VGND.n50 VGND.n49 0.0185556
R1523 VGND.n49 VGND.n48 0.0171667
R1524 VGND.n489 VGND.n1 0.0169949
R1525 VGND.n467 VGND.n466 0.0158374
R1526 VGND.n48 VGND.n47 0.0157778
R1527 VGND.n46 VGND.n45 0.013
R1528 VGND.n47 VGND.n46 0.013
R1529 VGND.n45 VGND.n44 0.0102222
R1530 VGND.n293 VGND.n281 0.00943
R1531 VGND.n115 VGND.n96 0.00911038
R1532 VGND.n44 VGND.n43 0.00874176
R1533 VGND.n445 VGND.n41 0.00816087
R1534 VGND.n43 VGND.n41 0.00744444
R1535 VGND.n424 VGND.n423 0.00285443
R1536 uo_out[0] uo_out[0].t1 984.356
R1537 uo_out[0].n0 uo_out[0].t2 582.378
R1538 uo_out[0].n1 uo_out[0].t3 566.953
R1539 uo_out[0].n8 uo_out[0].t0 478.87
R1540 uo_out[0].n1 uo_out[0].n0 424.161
R1541 uo_out[0].n3 uo_out[0].t4 294.557
R1542 uo_out[0].n3 uo_out[0].t5 211.01
R1543 uo_out[0].n2 uo_out[0].n0 204.481
R1544 uo_out[0] uo_out[0].n1 201.921
R1545 uo_out[0].n4 uo_out[0].n3 152
R1546 uo_out[0].n7 uo_out[0].n6 18.3079
R1547 uo_out[0].n5 uo_out[0].n4 17.6405
R1548 uo_out[0].n2 uo_out[0] 10.2405
R1549 uo_out[0] uo_out[0].n8 10.2405
R1550 uo_out[0].n8 uo_out[0].n7 7.5409
R1551 uo_out[0].n6 uo_out[0].n5 6.83545
R1552 uo_out[0].n7 uo_out[0].n2 5.01603
R1553 uo_out[0].n4 uo_out[0] 2.01193
R1554 uo_out[0].n6 uo_out[0] 1.31337
R1555 uo_out[0].n5 uo_out[0] 0.0793043
R1556 uo_out[1].n2 uo_out[1].t1 313.104
R1557 uo_out[1].n0 uo_out[1].t2 294.557
R1558 uo_out[1].t0 uo_out[1].n2 265.769
R1559 uo_out[1] uo_out[1].t0 262.318
R1560 uo_out[1].n0 uo_out[1].t3 211.01
R1561 uo_out[1].n1 uo_out[1].n0 152
R1562 uo_out[1].n5 uo_out[1] 12.6752
R1563 uo_out[1].n4 uo_out[1].n1 11.6411
R1564 uo_out[1].n4 uo_out[1].n3 9.3005
R1565 uo_out[1].n3 uo_out[1] 7.17626
R1566 uo_out[1].n3 uo_out[1].n2 4.84898
R1567 uo_out[1].n5 uo_out[1].n4 4.5029
R1568 uo_out[1].n1 uo_out[1] 1.37896
R1569 uo_out[1] uo_out[1].n5 0.0730806
R1570 uo_out[3].n0 uo_out[3].t1 313.104
R1571 uo_out[3].t0 uo_out[3].n0 265.769
R1572 uo_out[3] uo_out[3].t0 262.318
R1573 uo_out[3].n2 uo_out[3] 19.5328
R1574 uo_out[3].n2 uo_out[3].n1 13.8005
R1575 uo_out[3].n1 uo_out[3].n0 7.17626
R1576 uo_out[3].n1 uo_out[3] 4.84898
R1577 uo_out[3] uo_out[3].n2 0.0529194
C0 m1_10514_15880# m2_10514_15880# 0.104063p
C1 m2_12074_25760# m1_12074_25760# 0.152927p
C2 m3_12074_25760# m2_12074_25760# 98.466896f
C3 m3_10514_15880# m4_10514_15880# 65.3249f
C4 m3_12074_25760# m4_12074_25760# 95.99921f
C5 m3_10514_15880# m2_10514_15880# 67.004105f
C6 uo_out[0] VGND 9.161321f
C7 uo_out[3] VGND 2.06525f
C8 VDPWR VGND 0.167785p
C9 m4_10514_15880# VGND 11.0708f $ **FLOATING
C10 m4_12074_25760# VGND 8.74739f $ **FLOATING
C11 m3_10514_15880# VGND 12.571401f $ **FLOATING
C12 m3_12074_25760# VGND 10.2012f $ **FLOATING
C13 m2_10514_15880# VGND 11.5358f $ **FLOATING
C14 m2_12074_25760# VGND 9.56448f $ **FLOATING
C15 m1_10514_15880# VGND 32.9027f $ **FLOATING
C16 m1_12074_25760# VGND 40.2807f $ **FLOATING
C17 ring_0/skullfet_inverter_16.A VGND 4.53396f
C18 ring_0/skullfet_inverter_17.A VGND 4.70918f
C19 ring_0/skullfet_inverter_15.A VGND 4.82841f
C20 ring_0/skullfet_inverter_18.A VGND 4.90629f
C21 ring_0/skullfet_inverter_14.A VGND 4.98419f
C22 ring_0/skullfet_inverter_19.A VGND 4.923029f
C23 ring_0/skullfet_inverter_13.A VGND 4.78946f
C24 ring_0/skullfet_inverter_20.A VGND 4.72064f
C25 ring_0/skullfet_inverter_12.A VGND 5.60339f
C26 ring_0/skullfet_inverter_20.Y VGND 5.35745f
C27 ring_0/skullfet_inverter_11.A VGND 4.96291f
C28 ring_0/skullfet_inverter_1.A VGND 5.16765f
C29 ring_0/skullfet_inverter_10.A VGND 5.58737f
C30 ring_0/skullfet_inverter_2.A VGND 5.65285f
C31 ring_0/skullfet_inverter_9.A VGND 4.78733f
C32 ring_0/skullfet_inverter_3.A VGND 4.92041f
C33 ring_0/skullfet_inverter_4.A VGND 4.93544f
C34 ring_0/skullfet_inverter_8.A VGND 4.94116f
C35 ring_0/skullfet_inverter_7.A VGND 4.81796f
C36 ring_0/skullfet_inverter_6.A VGND 4.53217f
.ends

