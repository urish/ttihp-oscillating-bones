** sch_path: /home/uri/p/ttihp-oscillating-bones/xschem/testbench.sch
**.subckt testbench
x1 osc_out osc_div_2 osc_div_4 osc_div_8 tt_um_oscillating_bones
R21 VGND osc_out 1Meg m=1
R22 VGND osc_div_2 1Meg m=1
R23 VGND osc_div_4 1Meg m=1
R24 VGND osc_div_8 1Meg m=1
V2 0 VGND 0
V4 VDPWR VGND 1.2
**** begin user architecture code

.lib /home/uri/p/IHP-Open-PDK/ihp-sg13g2/libs.tech/ngspice/models/cornerMOSlv.lib mos_tt
.include /home/uri/p/IHP-Open-PDK/ihp-sg13g2/libs.ref/sg13g2_stdcell/spice/sg13g2_stdcell.spice



.param temp=27
.param mc_ok=1

.tran 50p 200n
.save all

.control
run

meas tran tdiff TRIG osc_out VAL=1.1 RISE=2 TARG osc_out VAL=1.1 RISE=3
let osc_freq_mhz = (1 / (tdiff) / 1e6)
save osc_freq_mhz

meas tran tdiff_div2 TRIG osc_div_2 VAL=1.1 RISE=2 TARG osc_div_2 VAL=1.1 RISE=3
let osc_div_2_freq_mhz = (1 / (tdiff_div2) / 1e6)
save osc_div_2_freq_mhz

meas tran tdiff_div4 TRIG osc_div_4 VAL=1.1 RISE=2 TARG osc_div_4 VAL=1.1 RISE=3
let osc_div_4_freq_mhz = (1 / (tdiff_div4) / 1e6)
save osc_div_4_freq_mhz

meas tran tdiff_div8 TRIG osc_div_8 VAL=1.1 RISE=2 TARG osc_div_8 VAL=1.1 RISE=3
let osc_div_8_freq_mhz = (1 / (tdiff_div8) / 1e6)
save osc_div_8_freq_mhz

write testbench.raw
.endc


**** end user architecture code
**.ends

* expanding   symbol:  tt_um_oscillating_bones.sym # of pins=4
** sym_path: /home/uri/p/ttihp-oscillating-bones/xschem/tt_um_oscillating_bones.sym
** sch_path: /home/uri/p/ttihp-oscillating-bones/xschem/tt_um_oscillating_bones.sch
.subckt tt_um_oscillating_bones uo_out[0] uo_out[1] uo_out[2] uo_out[3]
*.opin uo_out[1]
*.opin uo_out[0]
*.opin uo_out[2]
*.opin uo_out[3]
x22 uo_out[1] uo_out[2] uo_out[3] uo_out[0] VDPWR VGND freq_divider
x1 uo_out[0] ring
.ends


* expanding   symbol:  freq_divider.sym # of pins=6
** sym_path: /home/uri/p/ttihp-oscillating-bones/xschem/freq_divider.sym
** sch_path: /home/uri/p/ttihp-oscillating-bones/xschem/freq_divider.sch
.subckt freq_divider ODIV2 ODIV4 ODIV8 IN VDD VSS
*.ipin IN
*.opin ODIV2
*.opin ODIV4
*.opin ODIV8
*.ipin VDD
*.ipin VSS
x4 ODIV2 net3 IN net3 VDD VDD VSS sg13g2_dfrbp_2
x1 ODIV4 net1 ODIV2 net1 VDD VDD VSS sg13g2_dfrbp_2
x2 ODIV8 net2 ODIV4 net2 VDD VDD VSS sg13g2_dfrbp_2
.ends


* expanding   symbol:  ring.sym # of pins=1
** sym_path: /home/uri/p/ttihp-oscillating-bones/xschem/ring.sym
** sch_path: /home/uri/p/ttihp-oscillating-bones/xschem/ring.sch
.subckt ring ROSC_OUT
*.opin ROSC_OUT
x1 net20 net1 skullfet_inverter
x2 net1 net3 skullfet_inverter
x3 net3 net2 skullfet_inverter
x4 net2 ROSC_OUT skullfet_inverter
x5 ROSC_OUT net4 skullfet_inverter
x7 net5 net6 skullfet_inverter
x6 net4 net5 skullfet_inverter
x8 net6 net7 skullfet_inverter
x9 net7 net11 skullfet_inverter
x10 net11 net8 skullfet_inverter
x11 net8 net9 skullfet_inverter
x12 net9 net10 skullfet_inverter
x13 net10 net12 skullfet_inverter
x14 net12 net13 skullfet_inverter
x15 net13 net14 skullfet_inverter
x16 net14 net15 skullfet_inverter
x17 net15 net16 skullfet_inverter
x18 net16 net17 skullfet_inverter
x19 net17 net18 skullfet_inverter
x20 net18 net19 skullfet_inverter
x21 net19 net20 skullfet_inverter
**** begin user architecture code


* Set an initial condition on net1 (0.0001 V) to break symmetry and assist DC operating point convergence in ngspice
.ic V(net1)=0.0001


**** end user architecture code
.ends


* expanding   symbol:  skullfet_inverter.sym # of pins=2
** sym_path: /home/uri/p/ttihp-oscillating-bones/xschem/skullfet_inverter.sym
** sch_path: /home/uri/p/ttihp-oscillating-bones/xschem/skullfet_inverter.sch
.subckt skullfet_inverter A Y
*.ipin A
*.opin Y
XM1 Y A VDPWR VDPWR sg13_lv_pmos w=4.05u l=0.4u ng=1 m=1
XM2 Y A VGND VGND sg13_lv_nmos w=4.05u l=0.4u ng=1 m=1
.ends

.GLOBAL VGND
.GLOBAL VDPWR
.end
