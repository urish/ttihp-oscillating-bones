MACRO tt_um_oscillating_bones
  CLASS BLOCK ;
  FOREIGN tt_um_oscillating_bones ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 15.434999 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.429000 ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 5.000 5.000 6.500 220.760 ;
    END
  END VAPWR
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 3.000 5.000 4.500 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 2.500 220.760 ;
    END
  END VGND
  OBS
      LAYER nwell ;
        RECT 46.960 219.685 75.400 221.290 ;
      LAYER pwell ;
        RECT 47.155 219.165 49.920 219.395 ;
        RECT 51.460 219.165 52.370 219.385 ;
        RECT 47.155 218.485 55.885 219.165 ;
        RECT 55.905 218.570 56.335 219.355 ;
        RECT 56.365 218.570 56.795 219.355 ;
        RECT 56.815 219.165 59.580 219.395 ;
        RECT 61.120 219.165 62.030 219.385 ;
        RECT 56.815 218.485 65.545 219.165 ;
        RECT 65.565 218.570 65.995 219.355 ;
        RECT 66.025 218.570 66.455 219.355 ;
        RECT 66.475 219.165 69.240 219.395 ;
        RECT 70.780 219.165 71.690 219.385 ;
        RECT 66.475 218.485 75.205 219.165 ;
        RECT 55.575 218.295 55.745 218.485 ;
        RECT 65.235 218.295 65.405 218.485 ;
        RECT 74.895 218.295 75.065 218.485 ;
        RECT 37.570 208.740 43.290 214.520 ;
      LAYER nwell ;
        RECT 46.010 208.740 52.350 214.520 ;
      LAYER pwell ;
        RECT 46.830 162.360 52.610 168.080 ;
        RECT 61.250 168.020 67.030 173.740 ;
        RECT 76.700 169.180 82.480 174.900 ;
        RECT 34.710 152.690 40.490 158.410 ;
      LAYER nwell ;
        RECT 46.830 153.300 52.610 159.640 ;
        RECT 61.250 158.960 67.030 165.300 ;
        RECT 76.700 160.120 82.480 166.460 ;
      LAYER pwell ;
        RECT 91.810 165.730 97.590 171.450 ;
      LAYER nwell ;
        RECT 91.810 156.670 97.590 163.010 ;
      LAYER pwell ;
        RECT 105.240 157.980 111.020 163.700 ;
        RECT 25.970 141.890 31.750 147.610 ;
      LAYER nwell ;
        RECT 34.710 143.630 40.490 149.970 ;
        RECT 105.240 148.920 111.020 155.260 ;
      LAYER pwell ;
        RECT 115.780 146.620 121.560 152.340 ;
      LAYER nwell ;
        RECT 25.970 132.830 31.750 139.170 ;
        RECT 115.780 137.560 121.560 143.900 ;
      LAYER pwell ;
        RECT 122.960 131.250 128.740 136.970 ;
        RECT 21.410 125.080 27.190 130.800 ;
      LAYER nwell ;
        RECT 21.410 116.020 27.190 122.360 ;
        RECT 122.960 122.190 128.740 128.530 ;
      LAYER pwell ;
        RECT 126.820 114.330 132.600 120.050 ;
        RECT 17.410 108.580 23.190 114.300 ;
      LAYER nwell ;
        RECT 17.410 99.520 23.190 105.860 ;
        RECT 126.820 105.270 132.600 111.610 ;
      LAYER pwell ;
        RECT 22.930 91.770 28.710 97.490 ;
      LAYER nwell ;
        RECT 122.680 96.740 128.460 103.080 ;
        RECT 22.930 82.710 28.710 89.050 ;
        RECT 32.170 79.250 37.950 85.590 ;
        RECT 113.240 83.820 119.020 90.160 ;
      LAYER pwell ;
        RECT 122.680 88.300 128.460 94.020 ;
        RECT 32.170 70.810 37.950 76.530 ;
      LAYER nwell ;
        RECT 44.280 69.580 50.060 75.920 ;
        RECT 102.700 73.960 108.480 80.300 ;
      LAYER pwell ;
        RECT 113.240 75.380 119.020 81.100 ;
        RECT 44.280 61.140 50.060 66.860 ;
      LAYER nwell ;
        RECT 58.710 63.920 64.490 70.260 ;
        RECT 74.160 62.760 79.940 69.100 ;
        RECT 89.270 66.210 95.050 72.550 ;
      LAYER pwell ;
        RECT 102.700 65.520 108.480 71.240 ;
        RECT 58.710 55.480 64.490 61.200 ;
        RECT 74.160 54.320 79.940 60.040 ;
        RECT 89.270 57.770 95.050 63.490 ;
      LAYER li1 ;
        RECT 47.150 221.015 75.210 221.185 ;
        RECT 47.240 219.860 47.575 220.845 ;
        RECT 47.745 219.875 47.960 221.015 ;
        RECT 48.150 220.095 48.480 220.825 ;
        RECT 47.240 219.290 47.475 219.860 ;
        RECT 48.150 219.705 48.420 220.095 ;
        RECT 48.670 219.955 49.000 220.800 ;
        RECT 49.170 220.005 49.340 221.015 ;
        RECT 49.510 220.285 49.850 220.845 ;
        RECT 50.085 220.515 50.400 221.015 ;
        RECT 50.580 220.545 51.465 220.715 ;
        RECT 47.645 219.375 48.420 219.705 ;
        RECT 47.240 218.635 47.495 219.290 ;
        RECT 48.220 218.995 48.420 219.375 ;
        RECT 48.590 219.875 49.000 219.955 ;
        RECT 49.510 219.910 50.410 220.285 ;
        RECT 48.590 219.825 48.825 219.875 ;
        RECT 48.590 219.245 48.780 219.825 ;
        RECT 49.510 219.705 49.700 219.910 ;
        RECT 50.580 219.705 50.750 220.545 ;
        RECT 51.690 220.515 51.940 220.845 ;
        RECT 48.950 219.375 49.700 219.705 ;
        RECT 49.870 219.375 50.750 219.705 ;
        RECT 48.590 219.205 48.835 219.245 ;
        RECT 49.500 219.205 49.700 219.375 ;
        RECT 48.590 219.120 48.990 219.205 ;
        RECT 47.665 218.465 47.985 218.925 ;
        RECT 48.220 218.725 48.470 218.995 ;
        RECT 48.660 218.685 48.990 219.120 ;
        RECT 49.160 218.465 49.330 219.075 ;
        RECT 49.500 218.680 49.830 219.205 ;
        RECT 50.095 218.465 50.305 218.995 ;
        RECT 50.580 218.915 50.750 219.375 ;
        RECT 50.920 219.415 51.240 220.375 ;
        RECT 51.410 219.625 51.600 220.345 ;
        RECT 51.770 219.445 51.940 220.515 ;
        RECT 52.110 220.215 52.280 221.015 ;
        RECT 52.450 220.570 53.555 220.740 ;
        RECT 52.450 219.955 52.620 220.570 ;
        RECT 53.765 220.420 54.015 220.845 ;
        RECT 54.185 220.555 54.450 221.015 ;
        RECT 52.790 220.035 53.320 220.400 ;
        RECT 53.765 220.290 54.070 220.420 ;
        RECT 52.110 219.865 52.620 219.955 ;
        RECT 52.110 219.695 52.980 219.865 ;
        RECT 52.110 219.625 52.280 219.695 ;
        RECT 52.400 219.445 52.600 219.475 ;
        RECT 50.920 219.085 51.385 219.415 ;
        RECT 51.770 219.145 52.600 219.445 ;
        RECT 51.770 218.915 51.940 219.145 ;
        RECT 50.580 218.745 51.365 218.915 ;
        RECT 51.535 218.745 51.940 218.915 ;
        RECT 52.120 218.465 52.490 218.965 ;
        RECT 52.810 218.915 52.980 219.695 ;
        RECT 53.150 219.335 53.320 220.035 ;
        RECT 53.490 219.505 53.730 220.100 ;
        RECT 53.150 219.115 53.675 219.335 ;
        RECT 53.900 219.185 54.070 220.290 ;
        RECT 53.845 219.055 54.070 219.185 ;
        RECT 54.240 219.095 54.520 220.045 ;
        RECT 53.845 218.915 54.015 219.055 ;
        RECT 52.810 218.745 53.485 218.915 ;
        RECT 53.680 218.745 54.015 218.915 ;
        RECT 54.185 218.465 54.435 218.925 ;
        RECT 54.690 218.725 54.875 220.845 ;
        RECT 55.045 220.515 55.375 221.015 ;
        RECT 55.545 220.345 55.715 220.845 ;
        RECT 55.050 220.175 55.715 220.345 ;
        RECT 55.050 219.185 55.280 220.175 ;
        RECT 55.450 219.355 55.800 220.005 ;
        RECT 55.975 219.850 56.265 221.015 ;
        RECT 56.435 219.850 56.725 221.015 ;
        RECT 56.900 219.860 57.235 220.845 ;
        RECT 57.405 219.875 57.620 221.015 ;
        RECT 57.810 220.095 58.140 220.825 ;
        RECT 56.900 219.290 57.135 219.860 ;
        RECT 57.810 219.705 58.080 220.095 ;
        RECT 58.330 219.955 58.660 220.800 ;
        RECT 58.830 220.005 59.000 221.015 ;
        RECT 59.170 220.285 59.510 220.845 ;
        RECT 59.745 220.515 60.060 221.015 ;
        RECT 60.240 220.545 61.125 220.715 ;
        RECT 57.305 219.375 58.080 219.705 ;
        RECT 55.050 219.015 55.715 219.185 ;
        RECT 55.045 218.465 55.375 218.845 ;
        RECT 55.545 218.725 55.715 219.015 ;
        RECT 55.975 218.465 56.265 219.190 ;
        RECT 56.435 218.465 56.725 219.190 ;
        RECT 56.900 218.635 57.155 219.290 ;
        RECT 57.880 218.995 58.080 219.375 ;
        RECT 58.250 219.875 58.660 219.955 ;
        RECT 59.170 219.910 60.070 220.285 ;
        RECT 58.250 219.825 58.485 219.875 ;
        RECT 58.250 219.245 58.440 219.825 ;
        RECT 59.170 219.705 59.360 219.910 ;
        RECT 60.240 219.705 60.410 220.545 ;
        RECT 61.350 220.515 61.600 220.845 ;
        RECT 58.610 219.375 59.360 219.705 ;
        RECT 59.530 219.375 60.410 219.705 ;
        RECT 58.250 219.205 58.495 219.245 ;
        RECT 59.160 219.205 59.360 219.375 ;
        RECT 58.250 219.120 58.650 219.205 ;
        RECT 57.325 218.465 57.645 218.925 ;
        RECT 57.880 218.725 58.130 218.995 ;
        RECT 58.320 218.685 58.650 219.120 ;
        RECT 58.820 218.465 58.990 219.075 ;
        RECT 59.160 218.680 59.490 219.205 ;
        RECT 59.755 218.465 59.965 218.995 ;
        RECT 60.240 218.915 60.410 219.375 ;
        RECT 60.580 219.415 60.900 220.375 ;
        RECT 61.070 219.625 61.260 220.345 ;
        RECT 61.430 219.445 61.600 220.515 ;
        RECT 61.770 220.215 61.940 221.015 ;
        RECT 62.110 220.570 63.215 220.740 ;
        RECT 62.110 219.955 62.280 220.570 ;
        RECT 63.425 220.420 63.675 220.845 ;
        RECT 63.845 220.555 64.110 221.015 ;
        RECT 62.450 220.035 62.980 220.400 ;
        RECT 63.425 220.290 63.730 220.420 ;
        RECT 61.770 219.865 62.280 219.955 ;
        RECT 61.770 219.695 62.640 219.865 ;
        RECT 61.770 219.625 61.940 219.695 ;
        RECT 62.060 219.445 62.260 219.475 ;
        RECT 60.580 219.085 61.045 219.415 ;
        RECT 61.430 219.145 62.260 219.445 ;
        RECT 61.430 218.915 61.600 219.145 ;
        RECT 60.240 218.745 61.025 218.915 ;
        RECT 61.195 218.745 61.600 218.915 ;
        RECT 61.780 218.465 62.150 218.965 ;
        RECT 62.470 218.915 62.640 219.695 ;
        RECT 62.810 219.335 62.980 220.035 ;
        RECT 63.150 219.505 63.390 220.100 ;
        RECT 62.810 219.115 63.335 219.335 ;
        RECT 63.560 219.185 63.730 220.290 ;
        RECT 63.505 219.055 63.730 219.185 ;
        RECT 63.900 219.095 64.180 220.045 ;
        RECT 63.505 218.915 63.675 219.055 ;
        RECT 62.470 218.745 63.145 218.915 ;
        RECT 63.340 218.745 63.675 218.915 ;
        RECT 63.845 218.465 64.095 218.925 ;
        RECT 64.350 218.725 64.535 220.845 ;
        RECT 64.705 220.515 65.035 221.015 ;
        RECT 65.205 220.345 65.375 220.845 ;
        RECT 64.710 220.175 65.375 220.345 ;
        RECT 64.710 219.185 64.940 220.175 ;
        RECT 65.110 219.355 65.460 220.005 ;
        RECT 65.635 219.850 65.925 221.015 ;
        RECT 66.095 219.850 66.385 221.015 ;
        RECT 66.560 219.860 66.895 220.845 ;
        RECT 67.065 219.875 67.280 221.015 ;
        RECT 67.470 220.095 67.800 220.825 ;
        RECT 66.560 219.290 66.795 219.860 ;
        RECT 67.470 219.705 67.740 220.095 ;
        RECT 67.990 219.955 68.320 220.800 ;
        RECT 68.490 220.005 68.660 221.015 ;
        RECT 68.830 220.285 69.170 220.845 ;
        RECT 69.405 220.515 69.720 221.015 ;
        RECT 69.900 220.545 70.785 220.715 ;
        RECT 66.965 219.375 67.740 219.705 ;
        RECT 64.710 219.015 65.375 219.185 ;
        RECT 64.705 218.465 65.035 218.845 ;
        RECT 65.205 218.725 65.375 219.015 ;
        RECT 65.635 218.465 65.925 219.190 ;
        RECT 66.095 218.465 66.385 219.190 ;
        RECT 66.560 218.635 66.815 219.290 ;
        RECT 67.540 218.995 67.740 219.375 ;
        RECT 67.910 219.875 68.320 219.955 ;
        RECT 68.830 219.910 69.730 220.285 ;
        RECT 67.910 219.825 68.145 219.875 ;
        RECT 67.910 219.245 68.100 219.825 ;
        RECT 68.830 219.705 69.020 219.910 ;
        RECT 69.900 219.705 70.070 220.545 ;
        RECT 71.010 220.515 71.260 220.845 ;
        RECT 68.270 219.375 69.020 219.705 ;
        RECT 69.190 219.375 70.070 219.705 ;
        RECT 67.910 219.205 68.155 219.245 ;
        RECT 68.820 219.205 69.020 219.375 ;
        RECT 67.910 219.120 68.310 219.205 ;
        RECT 66.985 218.465 67.305 218.925 ;
        RECT 67.540 218.725 67.790 218.995 ;
        RECT 67.980 218.685 68.310 219.120 ;
        RECT 68.480 218.465 68.650 219.075 ;
        RECT 68.820 218.680 69.150 219.205 ;
        RECT 69.415 218.465 69.625 218.995 ;
        RECT 69.900 218.915 70.070 219.375 ;
        RECT 70.240 219.415 70.560 220.375 ;
        RECT 70.730 219.625 70.920 220.345 ;
        RECT 71.090 219.445 71.260 220.515 ;
        RECT 71.430 220.215 71.600 221.015 ;
        RECT 71.770 220.570 72.875 220.740 ;
        RECT 71.770 219.955 71.940 220.570 ;
        RECT 73.085 220.420 73.335 220.845 ;
        RECT 73.505 220.555 73.770 221.015 ;
        RECT 72.110 220.035 72.640 220.400 ;
        RECT 73.085 220.290 73.390 220.420 ;
        RECT 71.430 219.865 71.940 219.955 ;
        RECT 71.430 219.695 72.300 219.865 ;
        RECT 71.430 219.625 71.600 219.695 ;
        RECT 71.720 219.445 71.920 219.475 ;
        RECT 70.240 219.085 70.705 219.415 ;
        RECT 71.090 219.145 71.920 219.445 ;
        RECT 71.090 218.915 71.260 219.145 ;
        RECT 69.900 218.745 70.685 218.915 ;
        RECT 70.855 218.745 71.260 218.915 ;
        RECT 71.440 218.465 71.810 218.965 ;
        RECT 72.130 218.915 72.300 219.695 ;
        RECT 72.470 219.335 72.640 220.035 ;
        RECT 72.810 219.505 73.050 220.100 ;
        RECT 72.470 219.115 72.995 219.335 ;
        RECT 73.220 219.185 73.390 220.290 ;
        RECT 73.165 219.055 73.390 219.185 ;
        RECT 73.560 219.095 73.840 220.045 ;
        RECT 73.165 218.915 73.335 219.055 ;
        RECT 72.130 218.745 72.805 218.915 ;
        RECT 73.000 218.745 73.335 218.915 ;
        RECT 73.505 218.465 73.755 218.925 ;
        RECT 74.010 218.725 74.195 220.845 ;
        RECT 74.365 220.515 74.695 221.015 ;
        RECT 74.865 220.345 75.035 220.845 ;
        RECT 74.370 220.175 75.035 220.345 ;
        RECT 74.370 219.185 74.600 220.175 ;
        RECT 74.770 219.355 75.120 220.005 ;
        RECT 74.370 219.015 75.035 219.185 ;
        RECT 74.365 218.465 74.695 218.845 ;
        RECT 74.865 218.725 75.035 219.015 ;
        RECT 47.150 218.295 75.210 218.465 ;
        RECT 40.070 214.570 49.630 215.130 ;
        RECT 38.510 214.240 39.070 214.460 ;
        RECT 37.680 213.350 39.070 214.240 ;
        RECT 40.070 213.460 40.630 214.570 ;
        RECT 49.070 213.350 49.630 214.570 ;
        RECT 51.180 214.130 51.960 214.180 ;
        RECT 50.630 213.400 51.960 214.130 ;
        RECT 38.510 213.130 39.070 213.350 ;
        RECT 50.630 213.130 51.180 213.400 ;
        RECT 41.960 207.900 47.960 208.460 ;
        RECT 76.980 173.960 77.870 174.790 ;
        RECT 61.530 172.800 62.420 173.630 ;
        RECT 76.760 173.400 78.090 173.960 ;
        RECT 61.310 172.240 62.640 172.800 ;
        RECT 76.090 171.840 77.760 172.400 ;
        RECT 60.640 170.680 62.310 171.240 ;
        RECT 47.110 167.140 48.000 167.970 ;
        RECT 46.890 166.580 48.220 167.140 ;
        RECT 46.220 165.020 47.890 165.580 ;
        RECT 34.990 157.470 35.880 158.300 ;
        RECT 34.770 156.910 36.100 157.470 ;
        RECT 46.220 156.580 46.780 165.020 ;
        RECT 52.890 157.690 53.450 163.690 ;
        RECT 60.640 162.240 61.200 170.680 ;
        RECT 67.310 163.350 67.870 169.350 ;
        RECT 76.090 163.400 76.650 171.840 ;
        RECT 92.090 170.510 92.980 171.340 ;
        RECT 82.760 164.510 83.320 170.510 ;
        RECT 91.870 169.950 93.200 170.510 ;
        RECT 91.200 168.390 92.870 168.950 ;
        RECT 76.090 162.840 77.870 163.400 ;
        RECT 60.640 161.680 62.420 162.240 ;
        RECT 77.090 161.290 78.090 161.840 ;
        RECT 61.640 160.130 62.640 160.680 ;
        RECT 77.040 160.510 77.820 161.290 ;
        RECT 61.590 159.350 62.370 160.130 ;
        RECT 91.200 159.950 91.760 168.390 ;
        RECT 97.870 161.060 98.430 167.060 ;
        RECT 105.520 162.760 106.410 163.590 ;
        RECT 105.300 162.200 106.630 162.760 ;
        RECT 104.630 160.640 106.300 161.200 ;
        RECT 91.200 159.390 92.980 159.950 ;
        RECT 92.200 157.840 93.200 158.390 ;
        RECT 92.150 157.060 92.930 157.840 ;
        RECT 46.220 156.020 48.000 156.580 ;
        RECT 34.100 155.350 35.770 155.910 ;
        RECT 26.250 146.670 27.140 147.500 ;
        RECT 34.100 146.910 34.660 155.350 ;
        RECT 47.220 154.470 48.220 155.020 ;
        RECT 40.770 148.020 41.330 154.020 ;
        RECT 47.170 153.690 47.950 154.470 ;
        RECT 104.630 152.200 105.190 160.640 ;
        RECT 111.300 153.310 111.860 159.310 ;
        RECT 104.630 151.640 106.410 152.200 ;
        RECT 116.060 151.400 116.950 152.230 ;
        RECT 115.840 150.840 117.170 151.400 ;
        RECT 105.630 150.090 106.630 150.640 ;
        RECT 105.580 149.310 106.360 150.090 ;
        RECT 115.170 149.280 116.840 149.840 ;
        RECT 26.030 146.110 27.360 146.670 ;
        RECT 34.100 146.350 35.880 146.910 ;
        RECT 25.360 144.550 27.030 145.110 ;
        RECT 35.100 144.800 36.100 145.350 ;
        RECT 25.360 136.110 25.920 144.550 ;
        RECT 35.050 144.020 35.830 144.800 ;
        RECT 32.030 137.220 32.590 143.220 ;
        RECT 115.170 140.840 115.730 149.280 ;
        RECT 121.840 141.950 122.400 147.950 ;
        RECT 115.170 140.280 116.950 140.840 ;
        RECT 116.170 138.730 117.170 139.280 ;
        RECT 116.120 137.950 116.900 138.730 ;
        RECT 25.360 135.550 27.140 136.110 ;
        RECT 127.570 136.030 128.460 136.860 ;
        RECT 127.350 135.470 128.680 136.030 ;
        RECT 26.360 134.000 27.360 134.550 ;
        RECT 26.310 133.220 27.090 134.000 ;
        RECT 127.680 133.910 129.350 134.470 ;
        RECT 21.690 129.860 22.580 130.690 ;
        RECT 21.470 129.300 22.800 129.860 ;
        RECT 20.800 127.740 22.470 128.300 ;
        RECT 20.800 119.300 21.360 127.740 ;
        RECT 122.120 126.580 122.680 132.580 ;
        RECT 27.470 120.410 28.030 126.410 ;
        RECT 128.790 125.470 129.350 133.910 ;
        RECT 127.570 124.910 129.350 125.470 ;
        RECT 127.350 123.360 128.350 123.910 ;
        RECT 127.620 122.580 128.400 123.360 ;
        RECT 20.800 118.740 22.580 119.300 ;
        RECT 127.100 119.110 127.990 119.940 ;
        RECT 126.880 118.550 128.210 119.110 ;
        RECT 21.800 117.190 22.800 117.740 ;
        RECT 21.750 116.410 22.530 117.190 ;
        RECT 126.210 116.990 127.880 117.550 ;
        RECT 17.690 113.360 18.580 114.190 ;
        RECT 17.470 112.800 18.800 113.360 ;
        RECT 16.800 111.240 18.470 111.800 ;
        RECT 16.800 102.800 17.360 111.240 ;
        RECT 23.470 103.910 24.030 109.910 ;
        RECT 126.210 108.550 126.770 116.990 ;
        RECT 132.880 109.660 133.440 115.660 ;
        RECT 126.210 107.990 127.990 108.550 ;
        RECT 127.210 106.440 128.210 106.990 ;
        RECT 127.160 105.660 127.940 106.440 ;
        RECT 16.800 102.240 18.580 102.800 ;
        RECT 127.340 101.910 128.120 102.690 ;
        RECT 127.070 101.360 128.070 101.910 ;
        RECT 17.800 100.690 18.800 101.240 ;
        RECT 17.750 99.910 18.530 100.690 ;
        RECT 127.290 99.800 129.070 100.360 ;
        RECT 27.540 96.550 28.430 97.380 ;
        RECT 27.320 95.990 28.650 96.550 ;
        RECT 27.650 94.430 29.320 94.990 ;
        RECT 22.090 87.100 22.650 93.100 ;
        RECT 28.760 85.990 29.320 94.430 ;
        RECT 121.840 92.690 122.400 98.690 ;
        RECT 128.510 91.360 129.070 99.800 ;
        RECT 127.400 90.800 129.070 91.360 ;
        RECT 117.900 88.990 118.680 89.770 ;
        RECT 127.070 89.240 128.400 89.800 ;
        RECT 117.630 88.440 118.630 88.990 ;
        RECT 127.290 88.410 128.180 89.240 ;
        RECT 117.850 86.880 119.630 87.440 ;
        RECT 27.540 85.430 29.320 85.990 ;
        RECT 27.320 83.880 28.320 84.430 ;
        RECT 36.830 84.420 37.610 85.200 ;
        RECT 27.590 83.100 28.370 83.880 ;
        RECT 36.560 83.870 37.560 84.420 ;
        RECT 36.780 82.310 38.560 82.870 ;
        RECT 31.330 75.200 31.890 81.200 ;
        RECT 38.000 73.870 38.560 82.310 ;
        RECT 107.360 79.130 108.140 79.910 ;
        RECT 112.400 79.770 112.960 85.770 ;
        RECT 107.090 78.580 108.090 79.130 ;
        RECT 119.070 78.440 119.630 86.880 ;
        RECT 117.960 77.880 119.630 78.440 ;
        RECT 107.310 77.020 109.090 77.580 ;
        RECT 48.940 74.750 49.720 75.530 ;
        RECT 48.670 74.200 49.670 74.750 ;
        RECT 36.890 73.310 38.560 73.870 ;
        RECT 48.890 72.640 50.670 73.200 ;
        RECT 36.560 71.750 37.890 72.310 ;
        RECT 36.780 70.920 37.670 71.750 ;
        RECT 43.440 65.530 44.000 71.530 ;
        RECT 50.110 64.200 50.670 72.640 ;
        RECT 93.930 71.380 94.710 72.160 ;
        RECT 93.660 70.830 94.660 71.380 ;
        RECT 101.860 69.910 102.420 75.910 ;
        RECT 63.370 69.090 64.150 69.870 ;
        RECT 93.880 69.270 95.660 69.830 ;
        RECT 63.100 68.540 64.100 69.090 ;
        RECT 78.820 67.930 79.600 68.710 ;
        RECT 63.320 66.980 65.100 67.540 ;
        RECT 78.550 67.380 79.550 67.930 ;
        RECT 49.000 63.640 50.670 64.200 ;
        RECT 48.670 62.080 50.000 62.640 ;
        RECT 48.890 61.250 49.780 62.080 ;
        RECT 57.870 59.870 58.430 65.870 ;
        RECT 64.540 58.540 65.100 66.980 ;
        RECT 78.770 65.820 80.550 66.380 ;
        RECT 73.320 58.710 73.880 64.710 ;
        RECT 63.430 57.980 65.100 58.540 ;
        RECT 79.990 57.380 80.550 65.820 ;
        RECT 88.430 62.160 88.990 68.160 ;
        RECT 95.100 60.830 95.660 69.270 ;
        RECT 108.530 68.580 109.090 77.020 ;
        RECT 117.630 76.320 118.960 76.880 ;
        RECT 117.850 75.490 118.740 76.320 ;
        RECT 107.420 68.020 109.090 68.580 ;
        RECT 107.090 66.460 108.420 67.020 ;
        RECT 107.310 65.630 108.200 66.460 ;
        RECT 93.990 60.270 95.660 60.830 ;
        RECT 93.660 58.710 94.990 59.270 ;
        RECT 93.880 57.880 94.770 58.710 ;
        RECT 63.100 56.420 64.430 56.980 ;
        RECT 78.880 56.820 80.550 57.380 ;
        RECT 63.320 55.590 64.210 56.420 ;
        RECT 78.550 55.260 79.880 55.820 ;
        RECT 78.770 54.430 79.660 55.260 ;
      LAYER met1 ;
        RECT 74.895 221.340 76.660 221.345 ;
        RECT 47.150 220.865 76.660 221.340 ;
        RECT 47.150 220.860 75.210 220.865 ;
        RECT 51.360 220.320 51.650 220.365 ;
        RECT 52.930 220.320 53.220 220.365 ;
        RECT 55.030 220.320 55.320 220.365 ;
        RECT 51.360 220.180 55.320 220.320 ;
        RECT 51.360 220.135 51.650 220.180 ;
        RECT 52.930 220.135 53.220 220.180 ;
        RECT 55.030 220.135 55.320 220.180 ;
        RECT 61.020 220.320 61.310 220.365 ;
        RECT 62.590 220.320 62.880 220.365 ;
        RECT 64.690 220.320 64.980 220.365 ;
        RECT 61.020 220.180 64.980 220.320 ;
        RECT 61.020 220.135 61.310 220.180 ;
        RECT 62.590 220.135 62.880 220.180 ;
        RECT 64.690 220.135 64.980 220.180 ;
        RECT 70.680 220.320 70.970 220.365 ;
        RECT 72.250 220.320 72.540 220.365 ;
        RECT 74.350 220.320 74.640 220.365 ;
        RECT 70.680 220.180 74.640 220.320 ;
        RECT 70.680 220.135 70.970 220.180 ;
        RECT 72.250 220.135 72.540 220.180 ;
        RECT 74.350 220.135 74.640 220.180 ;
        RECT 47.240 219.870 47.530 220.100 ;
        RECT 50.925 219.980 51.215 220.025 ;
        RECT 53.445 219.980 53.735 220.025 ;
        RECT 54.635 219.980 54.925 220.025 ;
        RECT 47.350 219.640 47.490 219.870 ;
        RECT 50.925 219.840 54.925 219.980 ;
        RECT 56.895 219.870 57.185 220.100 ;
        RECT 60.585 219.980 60.875 220.025 ;
        RECT 63.105 219.980 63.395 220.025 ;
        RECT 64.295 219.980 64.585 220.025 ;
        RECT 50.925 219.795 51.215 219.840 ;
        RECT 53.445 219.795 53.735 219.840 ;
        RECT 54.635 219.795 54.925 219.840 ;
        RECT 54.210 219.640 54.500 219.680 ;
        RECT 47.350 219.500 54.500 219.640 ;
        RECT 54.210 219.450 54.500 219.500 ;
        RECT 55.500 219.425 55.790 219.655 ;
        RECT 57.005 219.640 57.145 219.870 ;
        RECT 60.585 219.840 64.585 219.980 ;
        RECT 66.560 219.870 66.850 220.100 ;
        RECT 70.245 219.980 70.535 220.025 ;
        RECT 72.765 219.980 73.055 220.025 ;
        RECT 73.955 219.980 74.245 220.025 ;
        RECT 60.585 219.795 60.875 219.840 ;
        RECT 63.105 219.795 63.395 219.840 ;
        RECT 64.295 219.795 64.585 219.840 ;
        RECT 63.865 219.640 64.155 219.680 ;
        RECT 57.005 219.500 64.155 219.640 ;
        RECT 63.865 219.450 64.155 219.500 ;
        RECT 65.160 219.425 65.450 219.655 ;
        RECT 66.670 219.640 66.810 219.870 ;
        RECT 70.245 219.840 74.245 219.980 ;
        RECT 74.800 219.840 75.080 219.900 ;
        RECT 70.245 219.795 70.535 219.840 ;
        RECT 72.765 219.795 73.055 219.840 ;
        RECT 73.955 219.795 74.245 219.840 ;
        RECT 73.530 219.640 73.820 219.680 ;
        RECT 66.670 219.500 73.820 219.640 ;
        RECT 73.530 219.450 73.820 219.500 ;
        RECT 74.740 219.455 75.100 219.840 ;
        RECT 48.620 218.770 49.050 219.090 ;
        RECT 55.560 219.075 55.730 219.425 ;
        RECT 58.335 219.075 58.625 219.105 ;
        RECT 55.560 219.020 58.625 219.075 ;
        RECT 65.220 219.075 65.390 219.425 ;
        RECT 74.800 219.395 75.080 219.455 ;
        RECT 67.940 219.075 68.350 219.120 ;
        RECT 55.560 218.905 58.710 219.020 ;
        RECT 65.220 218.905 68.350 219.075 ;
        RECT 58.300 218.760 58.710 218.905 ;
        RECT 67.940 218.860 68.350 218.905 ;
        RECT 45.790 218.140 75.210 218.620 ;
        RECT 51.520 216.130 52.180 216.690 ;
        RECT 44.410 215.630 45.060 215.725 ;
        RECT 36.510 214.685 37.110 215.185 ;
        RECT 38.400 214.680 39.010 215.130 ;
        RECT 38.510 214.020 39.010 214.680 ;
        RECT 43.040 214.450 43.640 214.750 ;
        RECT 44.240 214.570 45.240 215.630 ;
        RECT 45.740 214.450 46.640 214.750 ;
        RECT 50.740 214.570 51.350 215.130 ;
        RECT 39.140 213.550 40.940 213.850 ;
        RECT 42.740 213.550 43.940 214.450 ;
        RECT 45.440 214.150 46.940 214.450 ;
        RECT 45.440 213.850 46.640 214.150 ;
        RECT 45.440 213.550 46.340 213.850 ;
        RECT 48.740 213.550 50.540 213.850 ;
        RECT 50.740 213.740 51.180 214.570 ;
        RECT 38.540 213.250 41.840 213.550 ;
        RECT 43.040 213.250 44.240 213.550 ;
        RECT 38.540 212.950 40.640 213.250 ;
        RECT 41.240 212.950 41.840 213.250 ;
        RECT 43.640 212.950 44.240 213.250 ;
        RECT 45.440 212.950 46.040 213.550 ;
        RECT 47.840 213.250 51.140 213.550 ;
        RECT 47.840 212.950 48.440 213.250 ;
        RECT 49.040 212.950 51.140 213.250 ;
        RECT 38.240 212.650 40.340 212.950 ;
        RECT 37.940 212.050 40.340 212.650 ;
        RECT 41.540 212.650 42.140 212.950 ;
        RECT 43.640 212.650 44.540 212.950 ;
        RECT 41.540 212.350 43.040 212.650 ;
        RECT 43.940 212.350 44.540 212.650 ;
        RECT 45.140 212.350 45.740 212.950 ;
        RECT 47.540 212.650 48.140 212.950 ;
        RECT 46.640 212.350 48.140 212.650 ;
        RECT 49.340 212.650 51.440 212.950 ;
        RECT 41.240 212.050 42.740 212.350 ;
        RECT 37.940 211.750 41.840 212.050 ;
        RECT 42.140 211.750 43.040 212.050 ;
        RECT 44.240 211.750 45.440 212.350 ;
        RECT 46.940 212.050 48.440 212.350 ;
        RECT 49.340 212.050 51.740 212.650 ;
        RECT 46.640 211.750 47.540 212.050 ;
        RECT 47.840 211.750 51.740 212.050 ;
        RECT 37.940 211.450 41.540 211.750 ;
        RECT 42.140 211.450 42.740 211.750 ;
        RECT 44.540 211.450 45.140 211.750 ;
        RECT 46.940 211.450 47.540 211.750 ;
        RECT 48.140 211.450 51.740 211.750 ;
        RECT 37.940 211.150 41.840 211.450 ;
        RECT 42.140 211.150 43.040 211.450 ;
        RECT 37.940 210.250 40.340 211.150 ;
        RECT 41.240 210.850 42.740 211.150 ;
        RECT 44.240 210.850 45.440 211.450 ;
        RECT 46.640 211.150 47.540 211.450 ;
        RECT 47.840 211.150 51.740 211.450 ;
        RECT 46.940 210.850 48.440 211.150 ;
        RECT 41.540 210.550 43.040 210.850 ;
        RECT 43.940 210.550 44.540 210.850 ;
        RECT 41.540 210.250 42.140 210.550 ;
        RECT 38.540 209.950 40.640 210.250 ;
        RECT 41.240 209.950 42.140 210.250 ;
        RECT 43.640 210.250 44.540 210.550 ;
        RECT 45.140 210.250 45.740 210.850 ;
        RECT 46.640 210.550 48.140 210.850 ;
        RECT 47.540 210.250 48.140 210.550 ;
        RECT 49.340 210.250 51.740 211.150 ;
        RECT 43.640 209.950 44.240 210.250 ;
        RECT 38.540 209.650 41.540 209.950 ;
        RECT 43.040 209.650 44.240 209.950 ;
        RECT 45.440 209.650 46.040 210.250 ;
        RECT 47.540 209.950 48.440 210.250 ;
        RECT 49.040 209.950 51.140 210.250 ;
        RECT 48.140 209.650 51.140 209.950 ;
        RECT 39.140 209.350 40.940 209.650 ;
        RECT 42.740 208.750 43.940 209.650 ;
        RECT 45.440 209.350 46.340 209.650 ;
        RECT 48.740 209.350 50.540 209.650 ;
        RECT 45.440 209.050 46.640 209.350 ;
        RECT 45.440 208.750 46.940 209.050 ;
        RECT 43.040 208.450 43.640 208.750 ;
        RECT 44.240 207.350 45.240 208.460 ;
        RECT 45.440 208.450 46.640 208.750 ;
        RECT 44.480 161.140 44.980 207.350 ;
        RECT 78.570 174.230 80.970 174.530 ;
        RECT 76.090 173.960 76.540 174.070 ;
        RECT 76.090 173.460 77.200 173.960 ;
        RECT 78.270 173.930 80.970 174.230 ;
        RECT 63.120 173.070 65.520 173.370 ;
        RECT 77.670 173.330 81.570 173.930 ;
        RECT 60.640 172.800 61.090 172.910 ;
        RECT 60.640 172.300 61.750 172.800 ;
        RECT 62.820 172.770 65.520 173.070 ;
        RECT 62.220 172.170 66.120 172.770 ;
        RECT 61.920 170.970 66.420 172.170 ;
        RECT 77.370 172.130 81.870 173.330 ;
        RECT 77.370 171.830 78.270 172.130 ;
        RECT 77.370 171.530 77.970 171.830 ;
        RECT 61.920 170.670 62.820 170.970 ;
        RECT 61.920 170.370 62.520 170.670 ;
        RECT 62.220 170.070 62.520 170.370 ;
        RECT 63.720 170.070 64.620 170.970 ;
        RECT 65.520 170.670 66.420 170.970 ;
        RECT 65.820 170.370 66.420 170.670 ;
        RECT 77.670 171.230 77.970 171.530 ;
        RECT 79.170 171.230 80.070 172.130 ;
        RECT 80.970 171.830 81.870 172.130 ;
        RECT 81.270 171.530 81.870 171.830 ;
        RECT 81.270 171.230 81.570 171.530 ;
        RECT 77.670 170.930 78.270 171.230 ;
        RECT 78.870 170.930 80.370 171.230 ;
        RECT 80.970 170.930 81.570 171.230 ;
        RECT 77.670 170.630 79.470 170.930 ;
        RECT 79.770 170.630 81.270 170.930 ;
        RECT 93.680 170.780 96.080 171.080 ;
        RECT 65.820 170.070 66.120 170.370 ;
        RECT 78.270 170.330 79.170 170.630 ;
        RECT 80.070 170.330 81.270 170.630 ;
        RECT 91.200 170.510 91.650 170.620 ;
        RECT 62.220 169.770 62.820 170.070 ;
        RECT 63.420 169.770 64.920 170.070 ;
        RECT 65.520 169.770 66.120 170.070 ;
        RECT 62.220 169.470 64.020 169.770 ;
        RECT 64.320 169.470 65.820 169.770 ;
        RECT 78.570 169.730 80.670 170.330 ;
        RECT 91.200 170.010 92.310 170.510 ;
        RECT 93.380 170.480 96.080 170.780 ;
        RECT 92.780 169.880 96.680 170.480 ;
        RECT 62.820 169.170 63.720 169.470 ;
        RECT 64.620 169.170 65.820 169.470 ;
        RECT 76.770 169.430 77.670 169.730 ;
        RECT 78.570 169.430 78.870 169.730 ;
        RECT 79.170 169.430 79.470 169.730 ;
        RECT 79.770 169.430 80.070 169.730 ;
        RECT 80.370 169.430 80.670 169.730 ;
        RECT 81.570 169.430 82.470 169.730 ;
        RECT 63.120 168.570 65.220 169.170 ;
        RECT 76.470 168.830 77.970 169.430 ;
        RECT 81.270 168.830 82.770 169.430 ;
        RECT 61.320 168.270 62.220 168.570 ;
        RECT 63.120 168.270 63.420 168.570 ;
        RECT 63.720 168.270 64.020 168.570 ;
        RECT 64.320 168.270 64.620 168.570 ;
        RECT 64.920 168.270 65.220 168.570 ;
        RECT 66.120 168.270 67.020 168.570 ;
        RECT 76.770 168.530 78.570 168.830 ;
        RECT 80.670 168.530 82.470 168.830 ;
        RECT 92.480 168.680 96.980 169.880 ;
        RECT 48.700 167.410 51.100 167.710 ;
        RECT 61.020 167.670 62.520 168.270 ;
        RECT 65.820 167.670 67.320 168.270 ;
        RECT 77.670 168.230 78.870 168.530 ;
        RECT 80.370 168.230 81.570 168.530 ;
        RECT 92.480 168.380 93.380 168.680 ;
        RECT 75.590 167.960 76.650 168.230 ;
        RECT 46.220 167.140 46.670 167.250 ;
        RECT 46.220 166.640 47.330 167.140 ;
        RECT 48.400 167.110 51.100 167.410 ;
        RECT 61.320 167.370 63.120 167.670 ;
        RECT 65.220 167.370 67.020 167.670 ;
        RECT 71.510 167.460 76.650 167.960 ;
        RECT 78.270 167.930 79.470 168.230 ;
        RECT 79.770 167.930 80.970 168.230 ;
        RECT 82.760 167.960 83.870 168.230 ;
        RECT 92.480 168.080 93.080 168.380 ;
        RECT 47.800 166.510 51.700 167.110 ;
        RECT 62.220 167.070 63.420 167.370 ;
        RECT 64.920 167.070 66.120 167.370 ;
        RECT 60.140 166.800 61.200 167.070 ;
        RECT 47.500 165.310 52.000 166.510 ;
        RECT 47.500 165.010 48.400 165.310 ;
        RECT 47.500 164.710 48.100 165.010 ;
        RECT 47.800 164.410 48.100 164.710 ;
        RECT 49.300 164.410 50.200 165.310 ;
        RECT 51.100 165.010 52.000 165.310 ;
        RECT 51.400 164.710 52.000 165.010 ;
        RECT 56.750 166.300 61.200 166.800 ;
        RECT 62.820 166.770 64.020 167.070 ;
        RECT 64.320 166.770 65.520 167.070 ;
        RECT 67.310 166.800 68.420 167.070 ;
        RECT 67.310 166.780 68.810 166.800 ;
        RECT 71.510 166.780 72.010 167.460 ;
        RECT 75.590 167.230 76.650 167.460 ;
        RECT 78.870 167.330 80.370 167.930 ;
        RECT 82.760 167.460 87.420 167.960 ;
        RECT 78.270 167.030 79.470 167.330 ;
        RECT 79.770 167.030 80.970 167.330 ;
        RECT 82.760 167.230 83.870 167.460 ;
        RECT 51.400 164.410 51.700 164.710 ;
        RECT 47.800 164.110 48.400 164.410 ;
        RECT 49.000 164.110 50.500 164.410 ;
        RECT 51.100 164.110 51.700 164.410 ;
        RECT 47.800 163.810 49.600 164.110 ;
        RECT 49.900 163.810 51.400 164.110 ;
        RECT 48.400 163.510 49.300 163.810 ;
        RECT 50.200 163.510 51.400 163.810 ;
        RECT 48.700 162.910 50.800 163.510 ;
        RECT 46.900 162.610 47.800 162.910 ;
        RECT 48.700 162.610 49.000 162.910 ;
        RECT 49.300 162.610 49.600 162.910 ;
        RECT 49.900 162.610 50.200 162.910 ;
        RECT 50.500 162.610 50.800 162.910 ;
        RECT 51.700 162.610 52.600 162.910 ;
        RECT 46.600 162.010 48.100 162.610 ;
        RECT 51.400 162.010 52.900 162.610 ;
        RECT 46.900 161.710 48.700 162.010 ;
        RECT 50.800 161.710 52.600 162.010 ;
        RECT 47.800 161.410 49.000 161.710 ;
        RECT 50.500 161.410 51.700 161.710 ;
        RECT 45.720 161.140 46.780 161.410 ;
        RECT 43.590 160.640 46.780 161.140 ;
        RECT 48.400 161.110 49.600 161.410 ;
        RECT 49.900 161.110 51.100 161.410 ;
        RECT 52.890 161.160 54.000 161.410 ;
        RECT 56.750 161.160 57.250 166.300 ;
        RECT 60.140 166.070 61.200 166.300 ;
        RECT 63.420 166.170 64.920 166.770 ;
        RECT 67.310 166.280 72.010 166.780 ;
        RECT 76.770 166.730 78.870 167.030 ;
        RECT 80.370 166.730 82.770 167.030 ;
        RECT 76.470 166.430 78.270 166.730 ;
        RECT 80.970 166.430 82.770 166.730 ;
        RECT 62.820 165.870 64.020 166.170 ;
        RECT 64.320 165.870 65.520 166.170 ;
        RECT 67.310 166.070 68.420 166.280 ;
        RECT 76.470 166.130 77.670 166.430 ;
        RECT 81.570 166.130 82.770 166.430 ;
        RECT 61.320 165.570 63.420 165.870 ;
        RECT 64.920 165.570 67.320 165.870 ;
        RECT 76.470 165.830 77.370 166.130 ;
        RECT 81.870 165.830 82.770 166.130 ;
        RECT 61.020 165.270 62.820 165.570 ;
        RECT 65.520 165.270 67.320 165.570 ;
        RECT 76.770 165.530 77.070 165.830 ;
        RECT 78.570 165.530 78.870 165.830 ;
        RECT 79.170 165.530 79.470 165.830 ;
        RECT 79.770 165.530 80.070 165.830 ;
        RECT 80.370 165.530 80.670 165.830 ;
        RECT 82.170 165.530 82.470 165.830 ;
        RECT 61.020 164.970 62.220 165.270 ;
        RECT 66.120 164.970 67.320 165.270 ;
        RECT 61.020 164.670 61.920 164.970 ;
        RECT 66.420 164.670 67.320 164.970 ;
        RECT 78.570 164.930 80.670 165.530 ;
        RECT 61.320 164.370 61.620 164.670 ;
        RECT 63.120 164.370 63.420 164.670 ;
        RECT 63.720 164.370 64.020 164.670 ;
        RECT 64.320 164.370 64.620 164.670 ;
        RECT 64.920 164.370 65.220 164.670 ;
        RECT 66.720 164.370 67.020 164.670 ;
        RECT 78.270 164.630 79.170 164.930 ;
        RECT 80.070 164.630 81.270 164.930 ;
        RECT 63.120 163.770 65.220 164.370 ;
        RECT 77.670 164.330 79.470 164.630 ;
        RECT 79.770 164.330 81.270 164.630 ;
        RECT 86.920 164.510 87.420 167.460 ;
        RECT 92.780 167.780 93.080 168.080 ;
        RECT 94.280 167.780 95.180 168.680 ;
        RECT 96.080 168.380 96.980 168.680 ;
        RECT 96.380 168.080 96.980 168.380 ;
        RECT 96.380 167.780 96.680 168.080 ;
        RECT 92.780 167.480 93.380 167.780 ;
        RECT 93.980 167.480 95.480 167.780 ;
        RECT 96.080 167.480 96.680 167.780 ;
        RECT 92.780 167.180 94.580 167.480 ;
        RECT 94.880 167.180 96.380 167.480 ;
        RECT 93.380 166.880 94.280 167.180 ;
        RECT 95.180 166.880 96.380 167.180 ;
        RECT 93.680 166.280 95.780 166.880 ;
        RECT 91.880 165.980 92.780 166.280 ;
        RECT 93.680 165.980 93.980 166.280 ;
        RECT 94.280 165.980 94.580 166.280 ;
        RECT 94.880 165.980 95.180 166.280 ;
        RECT 95.480 165.980 95.780 166.280 ;
        RECT 96.680 165.980 97.580 166.280 ;
        RECT 91.580 165.380 93.080 165.980 ;
        RECT 96.380 165.380 97.880 165.980 ;
        RECT 91.880 165.080 93.680 165.380 ;
        RECT 95.780 165.080 97.580 165.380 ;
        RECT 92.780 164.780 93.980 165.080 ;
        RECT 95.480 164.780 96.680 165.080 ;
        RECT 90.700 164.510 91.760 164.780 ;
        RECT 77.670 164.030 78.270 164.330 ;
        RECT 78.870 164.030 80.370 164.330 ;
        RECT 80.970 164.030 81.570 164.330 ;
        RECT 62.820 163.470 63.720 163.770 ;
        RECT 64.620 163.470 65.820 163.770 ;
        RECT 77.670 163.730 77.970 164.030 ;
        RECT 62.220 163.170 64.020 163.470 ;
        RECT 64.320 163.170 65.820 163.470 ;
        RECT 77.370 163.430 77.970 163.730 ;
        RECT 62.220 162.870 62.820 163.170 ;
        RECT 63.420 162.870 64.920 163.170 ;
        RECT 65.520 162.870 66.120 163.170 ;
        RECT 62.220 162.570 62.520 162.870 ;
        RECT 36.580 157.740 38.980 158.040 ;
        RECT 34.100 157.470 34.550 157.580 ;
        RECT 34.100 156.970 35.210 157.470 ;
        RECT 36.280 157.440 38.980 157.740 ;
        RECT 35.680 156.840 39.580 157.440 ;
        RECT 35.380 155.640 39.880 156.840 ;
        RECT 35.380 155.340 36.280 155.640 ;
        RECT 35.380 155.040 35.980 155.340 ;
        RECT 35.680 154.740 35.980 155.040 ;
        RECT 37.180 154.740 38.080 155.640 ;
        RECT 38.980 155.340 39.880 155.640 ;
        RECT 39.280 155.040 39.880 155.340 ;
        RECT 39.280 154.740 39.580 155.040 ;
        RECT 35.680 154.440 36.280 154.740 ;
        RECT 36.880 154.440 38.380 154.740 ;
        RECT 38.980 154.440 39.580 154.740 ;
        RECT 35.680 154.140 37.480 154.440 ;
        RECT 37.780 154.140 39.280 154.440 ;
        RECT 36.280 153.840 37.180 154.140 ;
        RECT 38.080 153.840 39.280 154.140 ;
        RECT 36.580 153.240 38.680 153.840 ;
        RECT 34.780 152.940 35.680 153.240 ;
        RECT 36.580 152.940 36.880 153.240 ;
        RECT 37.180 152.940 37.480 153.240 ;
        RECT 37.780 152.940 38.080 153.240 ;
        RECT 38.380 152.940 38.680 153.240 ;
        RECT 39.580 152.940 40.480 153.240 ;
        RECT 34.480 152.340 35.980 152.940 ;
        RECT 39.280 152.340 40.780 152.940 ;
        RECT 34.780 152.040 36.580 152.340 ;
        RECT 38.680 152.040 40.480 152.340 ;
        RECT 35.680 151.740 36.880 152.040 ;
        RECT 38.380 151.740 39.580 152.040 ;
        RECT 33.600 151.470 34.660 151.740 ;
        RECT 33.100 150.740 34.660 151.470 ;
        RECT 36.280 151.440 37.480 151.740 ;
        RECT 37.780 151.440 38.980 151.740 ;
        RECT 40.770 151.480 41.880 151.740 ;
        RECT 43.590 151.480 44.090 160.640 ;
        RECT 45.720 160.410 46.780 160.640 ;
        RECT 49.000 160.510 50.500 161.110 ;
        RECT 52.890 160.660 57.250 161.160 ;
        RECT 61.920 162.270 62.520 162.570 ;
        RECT 61.920 161.970 62.820 162.270 ;
        RECT 63.720 161.970 64.620 162.870 ;
        RECT 65.820 162.570 66.120 162.870 ;
        RECT 77.370 163.130 78.270 163.430 ;
        RECT 79.170 163.130 80.070 164.030 ;
        RECT 81.270 163.730 81.570 164.030 ;
        RECT 86.920 164.010 91.760 164.510 ;
        RECT 93.380 164.480 94.580 164.780 ;
        RECT 94.880 164.480 96.080 164.780 ;
        RECT 97.870 164.510 98.980 164.780 ;
        RECT 90.700 163.780 91.760 164.010 ;
        RECT 93.980 163.880 95.480 164.480 ;
        RECT 97.870 164.010 101.510 164.510 ;
        RECT 81.270 163.430 81.870 163.730 ;
        RECT 93.380 163.580 94.580 163.880 ;
        RECT 94.880 163.580 96.080 163.880 ;
        RECT 97.870 163.780 98.980 164.010 ;
        RECT 80.970 163.130 81.870 163.430 ;
        RECT 91.880 163.280 93.980 163.580 ;
        RECT 95.480 163.280 97.880 163.580 ;
        RECT 65.820 162.270 66.420 162.570 ;
        RECT 65.520 161.970 66.420 162.270 ;
        RECT 61.920 160.770 66.420 161.970 ;
        RECT 77.370 161.930 81.870 163.130 ;
        RECT 91.580 162.980 93.380 163.280 ;
        RECT 96.080 162.980 97.880 163.280 ;
        RECT 91.580 162.680 92.780 162.980 ;
        RECT 96.680 162.680 97.880 162.980 ;
        RECT 91.580 162.380 92.480 162.680 ;
        RECT 96.980 162.380 97.880 162.680 ;
        RECT 91.880 162.080 92.180 162.380 ;
        RECT 93.680 162.080 93.980 162.380 ;
        RECT 94.280 162.080 94.580 162.380 ;
        RECT 94.880 162.080 95.180 162.380 ;
        RECT 95.480 162.080 95.780 162.380 ;
        RECT 97.280 162.080 97.580 162.380 ;
        RECT 76.090 161.290 77.480 161.730 ;
        RECT 77.670 161.330 81.570 161.930 ;
        RECT 93.680 161.480 95.780 162.080 ;
        RECT 76.090 161.120 76.650 161.290 ;
        RECT 78.270 161.030 80.970 161.330 ;
        RECT 93.380 161.180 94.280 161.480 ;
        RECT 95.180 161.180 96.380 161.480 ;
        RECT 52.890 160.640 54.390 160.660 ;
        RECT 48.400 160.210 49.600 160.510 ;
        RECT 49.900 160.210 51.100 160.510 ;
        RECT 52.890 160.410 54.000 160.640 ;
        RECT 46.900 159.910 49.000 160.210 ;
        RECT 50.500 159.910 52.900 160.210 ;
        RECT 60.640 160.130 62.030 160.570 ;
        RECT 62.220 160.170 66.120 160.770 ;
        RECT 78.570 160.730 80.970 161.030 ;
        RECT 92.780 160.880 94.580 161.180 ;
        RECT 94.880 160.880 96.380 161.180 ;
        RECT 92.780 160.580 93.380 160.880 ;
        RECT 93.980 160.580 95.480 160.880 ;
        RECT 96.080 160.580 96.680 160.880 ;
        RECT 92.780 160.280 93.080 160.580 ;
        RECT 60.640 159.960 61.200 160.130 ;
        RECT 46.600 159.610 48.400 159.910 ;
        RECT 51.100 159.610 52.900 159.910 ;
        RECT 62.820 159.870 65.520 160.170 ;
        RECT 46.600 159.310 47.800 159.610 ;
        RECT 51.700 159.310 52.900 159.610 ;
        RECT 63.120 159.570 65.520 159.870 ;
        RECT 92.480 159.980 93.080 160.280 ;
        RECT 92.480 159.680 93.380 159.980 ;
        RECT 94.280 159.680 95.180 160.580 ;
        RECT 96.380 160.280 96.680 160.580 ;
        RECT 96.380 159.980 96.980 160.280 ;
        RECT 96.080 159.680 96.980 159.980 ;
        RECT 46.600 159.010 47.500 159.310 ;
        RECT 52.000 159.010 52.900 159.310 ;
        RECT 46.900 158.710 47.200 159.010 ;
        RECT 48.700 158.710 49.000 159.010 ;
        RECT 49.300 158.710 49.600 159.010 ;
        RECT 49.900 158.710 50.200 159.010 ;
        RECT 50.500 158.710 50.800 159.010 ;
        RECT 52.300 158.710 52.600 159.010 ;
        RECT 48.700 158.110 50.800 158.710 ;
        RECT 92.480 158.480 96.980 159.680 ;
        RECT 48.400 157.810 49.300 158.110 ;
        RECT 50.200 157.810 51.400 158.110 ;
        RECT 47.800 157.510 49.600 157.810 ;
        RECT 49.900 157.510 51.400 157.810 ;
        RECT 91.200 157.840 92.590 158.280 ;
        RECT 92.780 157.880 96.680 158.480 ;
        RECT 91.200 157.670 91.760 157.840 ;
        RECT 93.380 157.580 96.080 157.880 ;
        RECT 47.800 157.210 48.400 157.510 ;
        RECT 49.000 157.210 50.500 157.510 ;
        RECT 51.100 157.210 51.700 157.510 ;
        RECT 93.680 157.280 96.080 157.580 ;
        RECT 47.800 156.910 48.100 157.210 ;
        RECT 47.500 156.610 48.100 156.910 ;
        RECT 47.500 156.310 48.400 156.610 ;
        RECT 49.300 156.310 50.200 157.210 ;
        RECT 51.400 156.910 51.700 157.210 ;
        RECT 51.400 156.610 52.000 156.910 ;
        RECT 51.100 156.310 52.000 156.610 ;
        RECT 47.500 155.110 52.000 156.310 ;
        RECT 101.010 156.750 101.510 164.010 ;
        RECT 107.110 163.030 109.510 163.330 ;
        RECT 104.630 162.760 105.080 162.870 ;
        RECT 104.630 162.260 105.740 162.760 ;
        RECT 106.810 162.730 109.510 163.030 ;
        RECT 106.210 162.130 110.110 162.730 ;
        RECT 105.910 160.930 110.410 162.130 ;
        RECT 105.910 160.630 106.810 160.930 ;
        RECT 105.910 160.330 106.510 160.630 ;
        RECT 106.210 160.030 106.510 160.330 ;
        RECT 107.710 160.030 108.610 160.930 ;
        RECT 109.510 160.630 110.410 160.930 ;
        RECT 109.810 160.330 110.410 160.630 ;
        RECT 109.810 160.030 110.110 160.330 ;
        RECT 106.210 159.730 106.810 160.030 ;
        RECT 107.410 159.730 108.910 160.030 ;
        RECT 109.510 159.730 110.110 160.030 ;
        RECT 106.210 159.430 108.010 159.730 ;
        RECT 108.310 159.430 109.810 159.730 ;
        RECT 106.810 159.130 107.710 159.430 ;
        RECT 108.610 159.130 109.810 159.430 ;
        RECT 107.110 158.530 109.210 159.130 ;
        RECT 105.310 158.230 106.210 158.530 ;
        RECT 107.110 158.230 107.410 158.530 ;
        RECT 107.710 158.230 108.010 158.530 ;
        RECT 108.310 158.230 108.610 158.530 ;
        RECT 108.910 158.230 109.210 158.530 ;
        RECT 110.110 158.230 111.010 158.530 ;
        RECT 105.010 157.630 106.510 158.230 ;
        RECT 109.810 157.630 111.310 158.230 ;
        RECT 105.310 157.330 107.110 157.630 ;
        RECT 109.210 157.330 111.010 157.630 ;
        RECT 106.210 157.030 107.410 157.330 ;
        RECT 108.910 157.030 110.110 157.330 ;
        RECT 104.130 156.760 105.190 157.030 ;
        RECT 103.630 156.750 105.190 156.760 ;
        RECT 101.010 156.260 105.190 156.750 ;
        RECT 106.810 156.730 108.010 157.030 ;
        RECT 108.310 156.730 109.510 157.030 ;
        RECT 111.300 156.760 112.410 157.030 ;
        RECT 101.010 156.250 103.970 156.260 ;
        RECT 104.130 156.030 105.190 156.260 ;
        RECT 107.410 156.130 108.910 156.730 ;
        RECT 111.300 156.260 113.520 156.760 ;
        RECT 106.810 155.830 108.010 156.130 ;
        RECT 108.310 155.830 109.510 156.130 ;
        RECT 111.300 156.030 112.410 156.260 ;
        RECT 105.310 155.530 107.410 155.830 ;
        RECT 108.910 155.530 111.310 155.830 ;
        RECT 105.010 155.230 106.810 155.530 ;
        RECT 109.510 155.230 111.310 155.530 ;
        RECT 46.220 154.470 47.610 154.910 ;
        RECT 47.800 154.510 51.700 155.110 ;
        RECT 105.010 154.930 106.210 155.230 ;
        RECT 110.110 154.930 111.310 155.230 ;
        RECT 105.010 154.630 105.910 154.930 ;
        RECT 110.410 154.630 111.310 154.930 ;
        RECT 46.220 154.300 46.780 154.470 ;
        RECT 48.400 154.210 51.100 154.510 ;
        RECT 105.310 154.330 105.610 154.630 ;
        RECT 107.110 154.330 107.410 154.630 ;
        RECT 107.710 154.330 108.010 154.630 ;
        RECT 108.310 154.330 108.610 154.630 ;
        RECT 108.910 154.330 109.210 154.630 ;
        RECT 110.710 154.330 111.010 154.630 ;
        RECT 48.700 153.910 51.100 154.210 ;
        RECT 107.110 153.730 109.210 154.330 ;
        RECT 106.810 153.430 107.710 153.730 ;
        RECT 108.610 153.430 109.810 153.730 ;
        RECT 106.210 153.130 108.010 153.430 ;
        RECT 108.310 153.130 109.810 153.430 ;
        RECT 106.210 152.830 106.810 153.130 ;
        RECT 107.410 152.830 108.910 153.130 ;
        RECT 109.510 152.830 110.110 153.130 ;
        RECT 106.210 152.530 106.510 152.830 ;
        RECT 36.880 150.840 38.380 151.440 ;
        RECT 40.770 150.980 44.090 151.480 ;
        RECT 105.910 152.230 106.510 152.530 ;
        RECT 105.910 151.930 106.810 152.230 ;
        RECT 107.710 151.930 108.610 152.830 ;
        RECT 109.810 152.530 110.110 152.830 ;
        RECT 109.810 152.230 110.410 152.530 ;
        RECT 109.510 151.930 110.410 152.230 ;
        RECT 40.770 150.970 42.270 150.980 ;
        RECT 27.840 146.940 30.240 147.240 ;
        RECT 25.360 146.670 25.810 146.780 ;
        RECT 25.360 146.170 26.470 146.670 ;
        RECT 27.540 146.640 30.240 146.940 ;
        RECT 26.940 146.040 30.840 146.640 ;
        RECT 26.640 144.840 31.140 146.040 ;
        RECT 26.640 144.540 27.540 144.840 ;
        RECT 26.640 144.240 27.240 144.540 ;
        RECT 26.940 143.940 27.240 144.240 ;
        RECT 28.440 143.940 29.340 144.840 ;
        RECT 30.240 144.540 31.140 144.840 ;
        RECT 30.540 144.240 31.140 144.540 ;
        RECT 30.540 143.940 30.840 144.240 ;
        RECT 26.940 143.640 27.540 143.940 ;
        RECT 28.140 143.640 29.640 143.940 ;
        RECT 30.240 143.640 30.840 143.940 ;
        RECT 26.940 143.340 28.740 143.640 ;
        RECT 29.040 143.340 30.540 143.640 ;
        RECT 27.540 143.040 28.440 143.340 ;
        RECT 29.340 143.040 30.540 143.340 ;
        RECT 27.840 142.440 29.940 143.040 ;
        RECT 26.040 142.140 26.940 142.440 ;
        RECT 27.840 142.140 28.140 142.440 ;
        RECT 28.440 142.140 28.740 142.440 ;
        RECT 29.040 142.140 29.340 142.440 ;
        RECT 29.640 142.140 29.940 142.440 ;
        RECT 30.840 142.140 31.740 142.440 ;
        RECT 25.740 141.540 27.240 142.140 ;
        RECT 30.540 141.540 32.040 142.140 ;
        RECT 26.040 141.240 27.840 141.540 ;
        RECT 29.940 141.240 31.740 141.540 ;
        RECT 26.940 140.940 28.140 141.240 ;
        RECT 29.640 140.940 30.840 141.240 ;
        RECT 33.100 140.940 33.600 150.740 ;
        RECT 36.280 150.540 37.480 150.840 ;
        RECT 37.780 150.540 38.980 150.840 ;
        RECT 40.770 150.740 41.880 150.970 ;
        RECT 105.910 150.730 110.410 151.930 ;
        RECT 34.780 150.240 36.880 150.540 ;
        RECT 38.380 150.240 40.780 150.540 ;
        RECT 34.480 149.940 36.280 150.240 ;
        RECT 38.980 149.940 40.780 150.240 ;
        RECT 34.480 149.640 35.680 149.940 ;
        RECT 39.580 149.640 40.780 149.940 ;
        RECT 34.480 149.340 35.380 149.640 ;
        RECT 39.880 149.340 40.780 149.640 ;
        RECT 34.780 149.040 35.080 149.340 ;
        RECT 36.580 149.040 36.880 149.340 ;
        RECT 37.180 149.040 37.480 149.340 ;
        RECT 37.780 149.040 38.080 149.340 ;
        RECT 38.380 149.040 38.680 149.340 ;
        RECT 40.180 149.040 40.480 149.340 ;
        RECT 36.580 148.440 38.680 149.040 ;
        RECT 36.280 148.140 37.180 148.440 ;
        RECT 38.080 148.140 39.280 148.440 ;
        RECT 66.380 148.410 84.060 150.620 ;
        RECT 104.630 150.090 106.020 150.530 ;
        RECT 106.210 150.130 110.110 150.730 ;
        RECT 104.630 149.920 105.190 150.090 ;
        RECT 106.810 149.830 109.510 150.130 ;
        RECT 107.110 149.530 109.510 149.830 ;
        RECT 35.680 147.840 37.480 148.140 ;
        RECT 37.780 147.840 39.280 148.140 ;
        RECT 35.680 147.540 36.280 147.840 ;
        RECT 36.880 147.540 38.380 147.840 ;
        RECT 38.980 147.540 39.580 147.840 ;
        RECT 35.680 147.240 35.980 147.540 ;
        RECT 35.380 146.940 35.980 147.240 ;
        RECT 35.380 146.640 36.280 146.940 ;
        RECT 37.180 146.640 38.080 147.540 ;
        RECT 39.280 147.240 39.580 147.540 ;
        RECT 39.280 146.940 39.880 147.240 ;
        RECT 38.980 146.640 39.880 146.940 ;
        RECT 35.380 145.440 39.880 146.640 ;
        RECT 64.170 146.200 84.060 148.410 ;
        RECT 34.100 144.800 35.490 145.240 ;
        RECT 35.680 144.840 39.580 145.440 ;
        RECT 34.100 144.630 34.660 144.800 ;
        RECT 36.280 144.540 38.980 144.840 ;
        RECT 36.580 144.240 38.980 144.540 ;
        RECT 59.750 141.780 88.480 146.200 ;
        RECT 113.020 145.400 113.520 156.260 ;
        RECT 117.650 151.670 120.050 151.970 ;
        RECT 115.170 151.400 115.620 151.510 ;
        RECT 115.170 150.900 116.280 151.400 ;
        RECT 117.350 151.370 120.050 151.670 ;
        RECT 116.750 150.770 120.650 151.370 ;
        RECT 116.450 149.570 120.950 150.770 ;
        RECT 116.450 149.270 117.350 149.570 ;
        RECT 116.450 148.970 117.050 149.270 ;
        RECT 116.750 148.670 117.050 148.970 ;
        RECT 118.250 148.670 119.150 149.570 ;
        RECT 120.050 149.270 120.950 149.570 ;
        RECT 120.350 148.970 120.950 149.270 ;
        RECT 120.350 148.670 120.650 148.970 ;
        RECT 116.750 148.370 117.350 148.670 ;
        RECT 117.950 148.370 119.450 148.670 ;
        RECT 120.050 148.370 120.650 148.670 ;
        RECT 116.750 148.070 118.550 148.370 ;
        RECT 118.850 148.070 120.350 148.370 ;
        RECT 117.350 147.770 118.250 148.070 ;
        RECT 119.150 147.770 120.350 148.070 ;
        RECT 117.650 147.170 119.750 147.770 ;
        RECT 115.850 146.870 116.750 147.170 ;
        RECT 117.650 146.870 117.950 147.170 ;
        RECT 118.250 146.870 118.550 147.170 ;
        RECT 118.850 146.870 119.150 147.170 ;
        RECT 119.450 146.870 119.750 147.170 ;
        RECT 120.650 146.870 121.550 147.170 ;
        RECT 115.550 146.270 117.050 146.870 ;
        RECT 120.350 146.270 121.850 146.870 ;
        RECT 115.850 145.970 117.650 146.270 ;
        RECT 119.750 145.970 121.550 146.270 ;
        RECT 116.750 145.670 117.950 145.970 ;
        RECT 119.450 145.670 120.650 145.970 ;
        RECT 114.670 145.400 115.730 145.670 ;
        RECT 113.020 144.900 115.730 145.400 ;
        RECT 117.350 145.370 118.550 145.670 ;
        RECT 118.850 145.370 120.050 145.670 ;
        RECT 121.840 145.400 122.950 145.670 ;
        RECT 114.670 144.670 115.730 144.900 ;
        RECT 117.950 144.770 119.450 145.370 ;
        RECT 121.840 144.900 124.180 145.400 ;
        RECT 117.350 144.470 118.550 144.770 ;
        RECT 118.850 144.470 120.050 144.770 ;
        RECT 121.840 144.670 122.950 144.900 ;
        RECT 115.850 144.170 117.950 144.470 ;
        RECT 119.450 144.170 121.850 144.470 ;
        RECT 115.550 143.870 117.350 144.170 ;
        RECT 120.050 143.870 121.850 144.170 ;
        RECT 115.550 143.570 116.750 143.870 ;
        RECT 120.650 143.570 121.850 143.870 ;
        RECT 115.550 143.270 116.450 143.570 ;
        RECT 120.950 143.270 121.850 143.570 ;
        RECT 115.850 142.970 116.150 143.270 ;
        RECT 117.650 142.970 117.950 143.270 ;
        RECT 118.250 142.970 118.550 143.270 ;
        RECT 118.850 142.970 119.150 143.270 ;
        RECT 119.450 142.970 119.750 143.270 ;
        RECT 121.250 142.970 121.550 143.270 ;
        RECT 117.650 142.370 119.750 142.970 ;
        RECT 117.350 142.070 118.250 142.370 ;
        RECT 119.150 142.070 120.350 142.370 ;
        RECT 24.860 140.670 25.920 140.940 ;
        RECT 24.360 139.940 25.920 140.670 ;
        RECT 27.540 140.640 28.740 140.940 ;
        RECT 29.040 140.640 30.240 140.940 ;
        RECT 28.140 140.040 29.640 140.640 ;
        RECT 32.030 140.210 33.600 140.940 ;
        RECT 32.030 140.170 33.530 140.210 ;
        RECT 24.360 131.860 24.860 139.940 ;
        RECT 27.540 139.740 28.740 140.040 ;
        RECT 29.040 139.740 30.240 140.040 ;
        RECT 32.030 139.940 33.140 140.170 ;
        RECT 26.040 139.440 28.140 139.740 ;
        RECT 29.640 139.440 32.040 139.740 ;
        RECT 25.740 139.140 27.540 139.440 ;
        RECT 30.240 139.140 32.040 139.440 ;
        RECT 25.740 138.840 26.940 139.140 ;
        RECT 30.840 138.840 32.040 139.140 ;
        RECT 25.740 138.540 26.640 138.840 ;
        RECT 31.140 138.540 32.040 138.840 ;
        RECT 26.040 138.240 26.340 138.540 ;
        RECT 27.840 138.240 28.140 138.540 ;
        RECT 28.440 138.240 28.740 138.540 ;
        RECT 29.040 138.240 29.340 138.540 ;
        RECT 29.640 138.240 29.940 138.540 ;
        RECT 31.440 138.240 31.740 138.540 ;
        RECT 27.840 137.640 29.940 138.240 ;
        RECT 27.540 137.340 28.440 137.640 ;
        RECT 29.340 137.340 30.540 137.640 ;
        RECT 26.940 137.040 28.740 137.340 ;
        RECT 29.040 137.040 30.540 137.340 ;
        RECT 26.940 136.740 27.540 137.040 ;
        RECT 28.140 136.740 29.640 137.040 ;
        RECT 30.240 136.740 30.840 137.040 ;
        RECT 26.940 136.440 27.240 136.740 ;
        RECT 26.640 136.140 27.240 136.440 ;
        RECT 26.640 135.840 27.540 136.140 ;
        RECT 28.440 135.840 29.340 136.740 ;
        RECT 30.540 136.440 30.840 136.740 ;
        RECT 30.540 136.140 31.140 136.440 ;
        RECT 30.240 135.840 31.140 136.140 ;
        RECT 26.640 134.640 31.140 135.840 ;
        RECT 25.360 134.000 26.750 134.440 ;
        RECT 26.940 134.040 30.840 134.640 ;
        RECT 25.360 133.830 25.920 134.000 ;
        RECT 27.540 133.740 30.240 134.040 ;
        RECT 27.840 133.440 30.240 133.740 ;
        RECT 57.540 132.940 90.690 141.780 ;
        RECT 116.750 141.770 118.550 142.070 ;
        RECT 118.850 141.770 120.350 142.070 ;
        RECT 116.750 141.470 117.350 141.770 ;
        RECT 117.950 141.470 119.450 141.770 ;
        RECT 120.050 141.470 120.650 141.770 ;
        RECT 116.750 141.170 117.050 141.470 ;
        RECT 116.450 140.870 117.050 141.170 ;
        RECT 116.450 140.570 117.350 140.870 ;
        RECT 118.250 140.570 119.150 141.470 ;
        RECT 120.350 141.170 120.650 141.470 ;
        RECT 120.350 140.870 120.950 141.170 ;
        RECT 120.050 140.570 120.950 140.870 ;
        RECT 116.450 139.370 120.950 140.570 ;
        RECT 115.170 138.730 116.560 139.170 ;
        RECT 116.750 138.770 120.650 139.370 ;
        RECT 115.170 138.560 115.730 138.730 ;
        RECT 117.350 138.470 120.050 138.770 ;
        RECT 117.650 138.170 120.050 138.470 ;
        RECT 123.680 138.670 124.180 144.900 ;
        RECT 123.680 138.170 130.340 138.670 ;
        RECT 124.470 136.300 126.870 136.600 ;
        RECT 124.470 136.000 127.170 136.300 ;
        RECT 128.900 136.030 129.350 136.140 ;
        RECT 123.870 135.400 127.770 136.000 ;
        RECT 128.240 135.530 129.350 136.030 ;
        RECT 123.570 134.200 128.070 135.400 ;
        RECT 123.570 133.900 124.470 134.200 ;
        RECT 123.570 133.600 124.170 133.900 ;
        RECT 123.870 133.300 124.170 133.600 ;
        RECT 125.370 133.300 126.270 134.200 ;
        RECT 127.170 133.900 128.070 134.200 ;
        RECT 127.470 133.600 128.070 133.900 ;
        RECT 127.470 133.300 127.770 133.600 ;
        RECT 123.870 133.000 124.470 133.300 ;
        RECT 125.070 133.000 126.570 133.300 ;
        RECT 127.170 133.000 127.770 133.300 ;
        RECT 24.360 131.360 28.910 131.860 ;
        RECT 23.280 130.130 25.680 130.430 ;
        RECT 20.800 129.860 21.250 129.970 ;
        RECT 20.800 129.360 21.910 129.860 ;
        RECT 22.980 129.830 25.680 130.130 ;
        RECT 22.380 129.230 26.280 129.830 ;
        RECT 22.080 128.030 26.580 129.230 ;
        RECT 22.080 127.730 22.980 128.030 ;
        RECT 22.080 127.430 22.680 127.730 ;
        RECT 22.380 127.130 22.680 127.430 ;
        RECT 23.880 127.130 24.780 128.030 ;
        RECT 25.680 127.730 26.580 128.030 ;
        RECT 25.980 127.430 26.580 127.730 ;
        RECT 25.980 127.130 26.280 127.430 ;
        RECT 22.380 126.830 22.980 127.130 ;
        RECT 23.580 126.830 25.080 127.130 ;
        RECT 25.680 126.830 26.280 127.130 ;
        RECT 22.380 126.530 24.180 126.830 ;
        RECT 24.480 126.530 25.980 126.830 ;
        RECT 22.980 126.230 23.880 126.530 ;
        RECT 24.780 126.230 25.980 126.530 ;
        RECT 23.280 125.630 25.380 126.230 ;
        RECT 21.480 125.330 22.380 125.630 ;
        RECT 23.280 125.330 23.580 125.630 ;
        RECT 23.880 125.330 24.180 125.630 ;
        RECT 24.480 125.330 24.780 125.630 ;
        RECT 25.080 125.330 25.380 125.630 ;
        RECT 26.280 125.330 27.180 125.630 ;
        RECT 21.180 124.730 22.680 125.330 ;
        RECT 25.980 124.730 27.480 125.330 ;
        RECT 21.480 124.430 23.280 124.730 ;
        RECT 25.380 124.430 27.180 124.730 ;
        RECT 22.380 124.130 23.580 124.430 ;
        RECT 25.080 124.130 26.280 124.430 ;
        RECT 28.410 124.130 28.910 131.360 ;
        RECT 57.540 130.730 64.170 132.940 ;
        RECT 57.540 128.520 61.960 130.730 ;
        RECT 19.470 123.860 19.970 123.930 ;
        RECT 20.300 123.860 21.360 124.130 ;
        RECT 19.470 123.360 21.360 123.860 ;
        RECT 22.980 123.830 24.180 124.130 ;
        RECT 24.480 123.830 25.680 124.130 ;
        RECT 27.470 123.860 28.910 124.130 ;
        RECT 59.750 126.310 61.960 128.520 ;
        RECT 70.800 126.310 77.430 132.940 ;
        RECT 84.060 130.730 90.690 132.940 ;
        RECT 124.170 132.700 125.670 133.000 ;
        RECT 125.970 132.700 127.770 133.000 ;
        RECT 124.170 132.400 125.370 132.700 ;
        RECT 126.270 132.400 127.170 132.700 ;
        RECT 124.770 131.800 126.870 132.400 ;
        RECT 122.970 131.500 123.870 131.800 ;
        RECT 124.770 131.500 125.070 131.800 ;
        RECT 125.370 131.500 125.670 131.800 ;
        RECT 125.970 131.500 126.270 131.800 ;
        RECT 126.570 131.500 126.870 131.800 ;
        RECT 127.770 131.500 128.670 131.800 ;
        RECT 122.670 130.900 124.170 131.500 ;
        RECT 127.470 130.900 128.970 131.500 ;
        RECT 86.270 128.520 90.690 130.730 ;
        RECT 122.970 130.600 124.770 130.900 ;
        RECT 126.870 130.600 128.670 130.900 ;
        RECT 123.870 130.300 125.070 130.600 ;
        RECT 126.570 130.300 127.770 130.600 ;
        RECT 129.840 130.300 130.340 138.170 ;
        RECT 121.570 130.030 122.680 130.300 ;
        RECT 121.180 129.300 122.680 130.030 ;
        RECT 124.470 130.000 125.670 130.300 ;
        RECT 125.970 130.000 127.170 130.300 ;
        RECT 128.790 130.030 130.340 130.300 ;
        RECT 125.070 129.400 126.570 130.000 ;
        RECT 128.790 129.530 130.350 130.030 ;
        RECT 86.270 126.310 88.480 128.520 ;
        RECT 59.750 124.100 64.170 126.310 ;
        RECT 68.590 124.100 79.640 126.310 ;
        RECT 84.060 124.100 88.480 126.310 ;
        RECT 19.470 114.940 19.970 123.360 ;
        RECT 20.300 123.130 21.360 123.360 ;
        RECT 23.580 123.230 25.080 123.830 ;
        RECT 27.470 123.360 28.970 123.860 ;
        RECT 22.980 122.930 24.180 123.230 ;
        RECT 24.480 122.930 25.680 123.230 ;
        RECT 27.470 123.130 28.580 123.360 ;
        RECT 21.480 122.630 23.580 122.930 ;
        RECT 25.080 122.630 27.480 122.930 ;
        RECT 21.180 122.330 22.980 122.630 ;
        RECT 25.680 122.330 27.480 122.630 ;
        RECT 21.180 122.030 22.380 122.330 ;
        RECT 26.280 122.030 27.480 122.330 ;
        RECT 21.180 121.730 22.080 122.030 ;
        RECT 26.580 121.730 27.480 122.030 ;
        RECT 59.750 121.890 73.010 124.100 ;
        RECT 75.220 121.890 86.270 124.100 ;
        RECT 21.480 121.430 21.780 121.730 ;
        RECT 23.280 121.430 23.580 121.730 ;
        RECT 23.880 121.430 24.180 121.730 ;
        RECT 24.480 121.430 24.780 121.730 ;
        RECT 25.080 121.430 25.380 121.730 ;
        RECT 26.880 121.430 27.180 121.730 ;
        RECT 23.280 120.830 25.380 121.430 ;
        RECT 22.980 120.530 23.880 120.830 ;
        RECT 24.780 120.530 25.980 120.830 ;
        RECT 22.380 120.230 24.180 120.530 ;
        RECT 24.480 120.230 25.980 120.530 ;
        RECT 22.380 119.930 22.980 120.230 ;
        RECT 23.580 119.930 25.080 120.230 ;
        RECT 25.680 119.930 26.280 120.230 ;
        RECT 22.380 119.630 22.680 119.930 ;
        RECT 22.080 119.330 22.680 119.630 ;
        RECT 22.080 119.030 22.980 119.330 ;
        RECT 23.880 119.030 24.780 119.930 ;
        RECT 25.980 119.630 26.280 119.930 ;
        RECT 64.170 119.680 70.800 121.890 ;
        RECT 77.430 119.680 86.270 121.890 ;
        RECT 25.980 119.330 26.580 119.630 ;
        RECT 25.680 119.030 26.580 119.330 ;
        RECT 22.080 117.830 26.580 119.030 ;
        RECT 20.800 117.190 22.190 117.630 ;
        RECT 22.380 117.230 26.280 117.830 ;
        RECT 20.800 117.020 21.360 117.190 ;
        RECT 22.980 116.930 25.680 117.230 ;
        RECT 23.280 116.630 25.680 116.930 ;
        RECT 66.380 115.260 81.850 119.680 ;
        RECT 19.470 114.440 24.970 114.940 ;
        RECT 7.470 112.910 9.070 114.410 ;
        RECT 19.280 113.630 21.680 113.930 ;
        RECT 16.800 113.360 17.250 113.470 ;
        RECT 16.800 112.860 17.910 113.360 ;
        RECT 18.980 113.330 21.680 113.630 ;
        RECT 18.380 112.730 22.280 113.330 ;
        RECT 18.080 111.530 22.580 112.730 ;
        RECT 18.080 111.230 18.980 111.530 ;
        RECT 18.080 110.930 18.680 111.230 ;
        RECT 18.380 110.630 18.680 110.930 ;
        RECT 19.880 110.630 20.780 111.530 ;
        RECT 21.680 111.230 22.580 111.530 ;
        RECT 21.980 110.930 22.580 111.230 ;
        RECT 21.980 110.630 22.280 110.930 ;
        RECT 18.380 110.330 18.980 110.630 ;
        RECT 19.580 110.330 21.080 110.630 ;
        RECT 21.680 110.330 22.280 110.630 ;
        RECT 18.380 110.030 20.180 110.330 ;
        RECT 20.480 110.030 21.980 110.330 ;
        RECT 18.980 109.730 19.880 110.030 ;
        RECT 20.780 109.730 21.980 110.030 ;
        RECT 19.280 109.130 21.380 109.730 ;
        RECT 17.480 108.830 18.380 109.130 ;
        RECT 19.280 108.830 19.580 109.130 ;
        RECT 19.880 108.830 20.180 109.130 ;
        RECT 20.480 108.830 20.780 109.130 ;
        RECT 21.080 108.830 21.380 109.130 ;
        RECT 22.280 108.830 23.180 109.130 ;
        RECT 17.180 108.230 18.680 108.830 ;
        RECT 21.980 108.230 23.480 108.830 ;
        RECT 17.480 107.930 19.280 108.230 ;
        RECT 21.380 107.930 23.180 108.230 ;
        RECT 18.380 107.630 19.580 107.930 ;
        RECT 21.080 107.630 22.280 107.930 ;
        RECT 24.470 107.630 24.970 114.440 ;
        RECT 53.120 113.050 59.750 115.260 ;
        RECT 66.380 113.050 68.590 115.260 ;
        RECT 70.800 113.050 73.010 115.260 ;
        RECT 75.220 113.050 77.430 115.260 ;
        RECT 79.640 113.050 81.850 115.260 ;
        RECT 88.480 113.050 95.110 115.260 ;
        RECT 121.180 113.110 121.680 129.300 ;
        RECT 124.470 129.100 125.670 129.400 ;
        RECT 125.970 129.100 127.170 129.400 ;
        RECT 128.790 129.300 129.850 129.530 ;
        RECT 122.670 128.800 125.070 129.100 ;
        RECT 126.570 128.800 128.670 129.100 ;
        RECT 122.670 128.500 124.470 128.800 ;
        RECT 127.170 128.500 128.970 128.800 ;
        RECT 122.670 128.200 123.870 128.500 ;
        RECT 127.770 128.200 128.970 128.500 ;
        RECT 122.670 127.900 123.570 128.200 ;
        RECT 128.070 127.900 128.970 128.200 ;
        RECT 122.970 127.600 123.270 127.900 ;
        RECT 124.770 127.600 125.070 127.900 ;
        RECT 125.370 127.600 125.670 127.900 ;
        RECT 125.970 127.600 126.270 127.900 ;
        RECT 126.570 127.600 126.870 127.900 ;
        RECT 128.370 127.600 128.670 127.900 ;
        RECT 124.770 127.000 126.870 127.600 ;
        RECT 124.170 126.700 125.370 127.000 ;
        RECT 126.270 126.700 127.170 127.000 ;
        RECT 124.170 126.400 125.670 126.700 ;
        RECT 125.970 126.400 127.770 126.700 ;
        RECT 123.870 126.100 124.470 126.400 ;
        RECT 125.070 126.100 126.570 126.400 ;
        RECT 127.170 126.100 127.770 126.400 ;
        RECT 123.870 125.800 124.170 126.100 ;
        RECT 123.570 125.500 124.170 125.800 ;
        RECT 123.570 125.200 124.470 125.500 ;
        RECT 125.370 125.200 126.270 126.100 ;
        RECT 127.470 125.800 127.770 126.100 ;
        RECT 127.470 125.500 128.070 125.800 ;
        RECT 127.170 125.200 128.070 125.500 ;
        RECT 123.570 124.000 128.070 125.200 ;
        RECT 123.870 123.400 127.770 124.000 ;
        RECT 124.470 123.100 127.170 123.400 ;
        RECT 127.960 123.360 129.350 123.800 ;
        RECT 128.790 123.190 129.350 123.360 ;
        RECT 124.470 122.800 126.870 123.100 ;
        RECT 128.690 119.380 131.090 119.680 ;
        RECT 126.210 119.110 126.660 119.220 ;
        RECT 126.210 118.610 127.320 119.110 ;
        RECT 128.390 119.080 131.090 119.380 ;
        RECT 127.790 118.480 131.690 119.080 ;
        RECT 127.490 117.280 131.990 118.480 ;
        RECT 127.490 116.980 128.390 117.280 ;
        RECT 127.490 116.680 128.090 116.980 ;
        RECT 127.790 116.380 128.090 116.680 ;
        RECT 129.290 116.380 130.190 117.280 ;
        RECT 131.090 116.980 131.990 117.280 ;
        RECT 131.390 116.680 131.990 116.980 ;
        RECT 131.390 116.380 131.690 116.680 ;
        RECT 127.790 116.080 128.390 116.380 ;
        RECT 128.990 116.080 130.490 116.380 ;
        RECT 131.090 116.080 131.690 116.380 ;
        RECT 127.790 115.780 129.590 116.080 ;
        RECT 129.890 115.780 131.390 116.080 ;
        RECT 128.390 115.480 129.290 115.780 ;
        RECT 130.190 115.480 131.390 115.780 ;
        RECT 128.690 114.880 130.790 115.480 ;
        RECT 126.890 114.580 127.790 114.880 ;
        RECT 128.690 114.580 128.990 114.880 ;
        RECT 129.290 114.580 129.590 114.880 ;
        RECT 129.890 114.580 130.190 114.880 ;
        RECT 130.490 114.580 130.790 114.880 ;
        RECT 131.690 114.580 132.590 114.880 ;
        RECT 126.590 113.980 128.090 114.580 ;
        RECT 131.390 113.980 132.890 114.580 ;
        RECT 126.890 113.680 128.690 113.980 ;
        RECT 130.790 113.680 132.590 113.980 ;
        RECT 127.790 113.380 128.990 113.680 ;
        RECT 130.490 113.380 131.690 113.680 ;
        RECT 125.710 113.110 126.770 113.380 ;
        RECT 50.910 108.630 61.960 113.050 ;
        RECT 86.270 108.630 97.320 113.050 ;
        RECT 121.180 112.610 126.770 113.110 ;
        RECT 128.390 113.080 129.590 113.380 ;
        RECT 129.890 113.080 131.090 113.380 ;
        RECT 132.880 113.110 133.990 113.380 ;
        RECT 125.710 112.380 126.770 112.610 ;
        RECT 128.990 112.480 130.490 113.080 ;
        RECT 132.880 112.610 135.290 113.110 ;
        RECT 128.390 112.180 129.590 112.480 ;
        RECT 129.890 112.180 131.090 112.480 ;
        RECT 132.880 112.380 133.990 112.610 ;
        RECT 126.890 111.880 128.990 112.180 ;
        RECT 130.490 111.880 132.890 112.180 ;
        RECT 126.590 111.580 128.390 111.880 ;
        RECT 131.090 111.580 132.890 111.880 ;
        RECT 126.590 111.280 127.790 111.580 ;
        RECT 131.690 111.280 132.890 111.580 ;
        RECT 126.590 110.980 127.490 111.280 ;
        RECT 131.990 110.980 132.890 111.280 ;
        RECT 126.890 110.680 127.190 110.980 ;
        RECT 128.690 110.680 128.990 110.980 ;
        RECT 129.290 110.680 129.590 110.980 ;
        RECT 129.890 110.680 130.190 110.980 ;
        RECT 130.490 110.680 130.790 110.980 ;
        RECT 132.290 110.680 132.590 110.980 ;
        RECT 128.690 110.080 130.790 110.680 ;
        RECT 128.390 109.780 129.290 110.080 ;
        RECT 130.190 109.780 131.390 110.080 ;
        RECT 127.790 109.480 129.590 109.780 ;
        RECT 129.890 109.480 131.390 109.780 ;
        RECT 127.790 109.180 128.390 109.480 ;
        RECT 128.990 109.180 130.490 109.480 ;
        RECT 131.090 109.180 131.690 109.480 ;
        RECT 127.790 108.880 128.090 109.180 ;
        RECT 16.300 107.360 17.360 107.630 ;
        RECT 15.800 106.630 17.360 107.360 ;
        RECT 18.980 107.330 20.180 107.630 ;
        RECT 20.480 107.330 21.680 107.630 ;
        RECT 19.580 106.730 21.080 107.330 ;
        RECT 23.470 106.860 24.970 107.630 ;
        RECT 15.800 97.460 16.300 106.630 ;
        RECT 18.980 106.430 20.180 106.730 ;
        RECT 20.480 106.430 21.680 106.730 ;
        RECT 23.470 106.630 24.580 106.860 ;
        RECT 17.480 106.130 19.580 106.430 ;
        RECT 21.080 106.130 23.480 106.430 ;
        RECT 53.120 106.420 66.380 108.630 ;
        RECT 81.850 106.420 95.110 108.630 ;
        RECT 127.490 108.580 128.090 108.880 ;
        RECT 127.490 108.280 128.390 108.580 ;
        RECT 129.290 108.280 130.190 109.180 ;
        RECT 131.390 108.880 131.690 109.180 ;
        RECT 131.390 108.580 131.990 108.880 ;
        RECT 131.090 108.280 131.990 108.580 ;
        RECT 127.490 107.080 131.990 108.280 ;
        RECT 126.210 106.440 127.600 106.880 ;
        RECT 127.790 106.480 131.690 107.080 ;
        RECT 17.180 105.830 18.980 106.130 ;
        RECT 21.680 105.830 23.480 106.130 ;
        RECT 17.180 105.530 18.380 105.830 ;
        RECT 22.280 105.530 23.480 105.830 ;
        RECT 17.180 105.230 18.080 105.530 ;
        RECT 22.580 105.230 23.480 105.530 ;
        RECT 17.480 104.930 17.780 105.230 ;
        RECT 19.280 104.930 19.580 105.230 ;
        RECT 19.880 104.930 20.180 105.230 ;
        RECT 20.480 104.930 20.780 105.230 ;
        RECT 21.080 104.930 21.380 105.230 ;
        RECT 22.880 104.930 23.180 105.230 ;
        RECT 19.280 104.330 21.380 104.930 ;
        RECT 18.980 104.030 19.880 104.330 ;
        RECT 20.780 104.030 21.980 104.330 ;
        RECT 59.750 104.210 68.590 106.420 ;
        RECT 79.640 104.210 88.480 106.420 ;
        RECT 126.210 106.270 126.770 106.440 ;
        RECT 128.390 106.180 131.090 106.480 ;
        RECT 128.690 105.880 131.090 106.180 ;
        RECT 134.790 104.710 135.290 112.610 ;
        RECT 129.520 104.210 135.290 104.710 ;
        RECT 18.380 103.730 20.180 104.030 ;
        RECT 20.480 103.730 21.980 104.030 ;
        RECT 18.380 103.430 18.980 103.730 ;
        RECT 19.580 103.430 21.080 103.730 ;
        RECT 21.680 103.430 22.280 103.730 ;
        RECT 18.380 103.130 18.680 103.430 ;
        RECT 18.080 102.830 18.680 103.130 ;
        RECT 18.080 102.530 18.980 102.830 ;
        RECT 19.880 102.530 20.780 103.430 ;
        RECT 21.980 103.130 22.280 103.430 ;
        RECT 21.980 102.830 22.580 103.130 ;
        RECT 21.680 102.530 22.580 102.830 ;
        RECT 18.080 101.330 22.580 102.530 ;
        RECT 64.170 102.000 73.010 104.210 ;
        RECT 75.220 102.000 84.060 104.210 ;
        RECT 124.190 102.170 126.590 102.470 ;
        RECT 16.800 100.690 18.190 101.130 ;
        RECT 18.380 100.730 22.280 101.330 ;
        RECT 16.800 100.520 17.360 100.690 ;
        RECT 18.980 100.430 21.680 100.730 ;
        RECT 19.280 100.130 21.680 100.430 ;
        RECT 68.590 97.580 79.640 102.000 ;
        RECT 124.190 101.870 126.890 102.170 ;
        RECT 128.510 101.910 129.070 102.080 ;
        RECT 123.590 101.270 127.490 101.870 ;
        RECT 127.680 101.470 129.070 101.910 ;
        RECT 123.290 100.070 127.790 101.270 ;
        RECT 123.290 99.770 124.190 100.070 ;
        RECT 123.290 99.470 123.890 99.770 ;
        RECT 123.590 99.170 123.890 99.470 ;
        RECT 125.090 99.170 125.990 100.070 ;
        RECT 126.890 99.770 127.790 100.070 ;
        RECT 127.190 99.470 127.790 99.770 ;
        RECT 127.190 99.170 127.490 99.470 ;
        RECT 123.590 98.870 124.190 99.170 ;
        RECT 124.790 98.870 126.290 99.170 ;
        RECT 126.890 98.870 127.490 99.170 ;
        RECT 123.890 98.570 125.390 98.870 ;
        RECT 125.690 98.570 127.490 98.870 ;
        RECT 123.890 98.270 125.090 98.570 ;
        RECT 125.990 98.270 126.890 98.570 ;
        RECT 124.490 97.670 126.590 98.270 ;
        RECT 15.800 96.960 19.830 97.460 ;
        RECT 19.330 90.590 19.830 96.960 ;
        RECT 24.440 96.820 26.840 97.120 ;
        RECT 24.440 96.520 27.140 96.820 ;
        RECT 28.870 96.550 29.320 96.660 ;
        RECT 23.840 95.920 27.740 96.520 ;
        RECT 28.210 96.050 29.320 96.550 ;
        RECT 23.540 94.720 28.040 95.920 ;
        RECT 64.170 95.370 73.010 97.580 ;
        RECT 75.220 95.370 84.060 97.580 ;
        RECT 122.690 97.370 122.990 97.670 ;
        RECT 124.490 97.370 124.790 97.670 ;
        RECT 125.090 97.370 125.390 97.670 ;
        RECT 125.690 97.370 125.990 97.670 ;
        RECT 126.290 97.370 126.590 97.670 ;
        RECT 128.090 97.370 128.390 97.670 ;
        RECT 122.390 97.070 123.290 97.370 ;
        RECT 127.790 97.070 128.690 97.370 ;
        RECT 122.390 96.770 123.590 97.070 ;
        RECT 127.490 96.770 128.690 97.070 ;
        RECT 122.390 96.470 124.190 96.770 ;
        RECT 126.890 96.470 128.690 96.770 ;
        RECT 122.390 96.170 124.790 96.470 ;
        RECT 126.290 96.170 128.390 96.470 ;
        RECT 121.290 95.790 122.400 95.970 ;
        RECT 124.190 95.870 125.390 96.170 ;
        RECT 125.690 95.870 126.890 96.170 ;
        RECT 129.520 95.970 130.020 104.210 ;
        RECT 23.540 94.420 24.440 94.720 ;
        RECT 23.540 94.120 24.140 94.420 ;
        RECT 23.840 93.820 24.140 94.120 ;
        RECT 25.340 93.820 26.240 94.720 ;
        RECT 27.140 94.420 28.040 94.720 ;
        RECT 27.440 94.120 28.040 94.420 ;
        RECT 27.440 93.820 27.740 94.120 ;
        RECT 23.840 93.520 24.440 93.820 ;
        RECT 25.040 93.520 26.540 93.820 ;
        RECT 27.140 93.520 27.740 93.820 ;
        RECT 24.140 93.220 25.640 93.520 ;
        RECT 25.940 93.220 27.740 93.520 ;
        RECT 24.140 92.920 25.340 93.220 ;
        RECT 26.240 92.920 27.140 93.220 ;
        RECT 53.120 93.160 68.590 95.370 ;
        RECT 79.640 93.160 97.320 95.370 ;
        RECT 24.740 92.320 26.840 92.920 ;
        RECT 22.940 92.020 23.840 92.320 ;
        RECT 24.740 92.020 25.040 92.320 ;
        RECT 25.340 92.020 25.640 92.320 ;
        RECT 25.940 92.020 26.240 92.320 ;
        RECT 26.540 92.020 26.840 92.320 ;
        RECT 27.740 92.020 28.640 92.320 ;
        RECT 22.640 91.420 24.140 92.020 ;
        RECT 27.440 91.420 28.940 92.020 ;
        RECT 22.940 91.120 24.740 91.420 ;
        RECT 26.840 91.120 28.640 91.420 ;
        RECT 23.840 90.820 25.040 91.120 ;
        RECT 26.540 90.820 27.740 91.120 ;
        RECT 50.910 90.950 64.170 93.160 ;
        RECT 84.060 90.950 97.320 93.160 ;
        RECT 21.540 90.590 22.650 90.820 ;
        RECT 19.330 90.090 22.650 90.590 ;
        RECT 24.440 90.520 25.640 90.820 ;
        RECT 25.940 90.520 27.140 90.820 ;
        RECT 21.540 89.820 22.650 90.090 ;
        RECT 25.040 89.920 26.540 90.520 ;
        RECT 28.760 90.490 29.820 90.820 ;
        RECT 28.760 89.990 30.780 90.490 ;
        RECT 24.440 89.620 25.640 89.920 ;
        RECT 25.940 89.620 27.140 89.920 ;
        RECT 28.760 89.820 29.820 89.990 ;
        RECT 22.640 89.320 25.040 89.620 ;
        RECT 26.540 89.320 28.640 89.620 ;
        RECT 22.640 89.020 24.440 89.320 ;
        RECT 27.140 89.020 28.940 89.320 ;
        RECT 22.640 88.720 23.840 89.020 ;
        RECT 27.740 88.720 28.940 89.020 ;
        RECT 22.640 88.420 23.540 88.720 ;
        RECT 28.040 88.420 28.940 88.720 ;
        RECT 22.940 88.120 23.240 88.420 ;
        RECT 24.740 88.120 25.040 88.420 ;
        RECT 25.340 88.120 25.640 88.420 ;
        RECT 25.940 88.120 26.240 88.420 ;
        RECT 26.540 88.120 26.840 88.420 ;
        RECT 28.340 88.120 28.640 88.420 ;
        RECT 24.740 87.520 26.840 88.120 ;
        RECT 24.140 87.220 25.340 87.520 ;
        RECT 26.240 87.220 27.140 87.520 ;
        RECT 24.140 86.920 25.640 87.220 ;
        RECT 25.940 86.920 27.740 87.220 ;
        RECT 23.840 86.620 24.440 86.920 ;
        RECT 25.040 86.620 26.540 86.920 ;
        RECT 27.140 86.620 27.740 86.920 ;
        RECT 23.840 86.320 24.140 86.620 ;
        RECT 23.540 86.020 24.140 86.320 ;
        RECT 23.540 85.720 24.440 86.020 ;
        RECT 25.340 85.720 26.240 86.620 ;
        RECT 27.440 86.320 27.740 86.620 ;
        RECT 27.440 86.020 28.040 86.320 ;
        RECT 27.140 85.720 28.040 86.020 ;
        RECT 23.540 84.520 28.040 85.720 ;
        RECT 23.840 83.920 27.740 84.520 ;
        RECT 24.440 83.620 27.140 83.920 ;
        RECT 27.930 83.880 29.320 84.320 ;
        RECT 28.760 83.710 29.320 83.880 ;
        RECT 24.440 83.320 26.840 83.620 ;
        RECT 30.280 78.480 30.780 89.990 ;
        RECT 50.910 88.740 59.750 90.950 ;
        RECT 88.480 88.740 97.320 90.950 ;
        RECT 120.420 95.290 122.400 95.790 ;
        RECT 114.750 89.250 117.150 89.550 ;
        RECT 114.750 88.950 117.450 89.250 ;
        RECT 119.070 88.990 119.630 89.160 ;
        RECT 50.910 86.530 57.540 88.740 ;
        RECT 90.690 86.530 97.320 88.740 ;
        RECT 114.150 88.350 118.050 88.950 ;
        RECT 118.240 88.550 119.630 88.990 ;
        RECT 113.850 87.150 118.350 88.350 ;
        RECT 113.850 86.850 114.750 87.150 ;
        RECT 113.850 86.550 114.450 86.850 ;
        RECT 33.680 84.680 36.080 84.980 ;
        RECT 33.680 84.380 36.380 84.680 ;
        RECT 38.000 84.420 38.560 84.590 ;
        RECT 33.080 83.780 36.980 84.380 ;
        RECT 37.170 83.980 38.560 84.420 ;
        RECT 53.120 84.320 55.330 86.530 ;
        RECT 92.900 84.320 95.110 86.530 ;
        RECT 114.150 86.250 114.450 86.550 ;
        RECT 115.650 86.250 116.550 87.150 ;
        RECT 117.450 86.850 118.350 87.150 ;
        RECT 117.750 86.550 118.350 86.850 ;
        RECT 117.750 86.250 118.050 86.550 ;
        RECT 114.150 85.950 114.750 86.250 ;
        RECT 115.350 85.950 116.850 86.250 ;
        RECT 117.450 85.950 118.050 86.250 ;
        RECT 114.450 85.650 115.950 85.950 ;
        RECT 116.250 85.650 118.050 85.950 ;
        RECT 114.450 85.350 115.650 85.650 ;
        RECT 116.550 85.350 117.450 85.650 ;
        RECT 115.050 84.750 117.150 85.350 ;
        RECT 113.250 84.450 113.550 84.750 ;
        RECT 115.050 84.450 115.350 84.750 ;
        RECT 115.650 84.450 115.950 84.750 ;
        RECT 116.250 84.450 116.550 84.750 ;
        RECT 116.850 84.450 117.150 84.750 ;
        RECT 118.650 84.450 118.950 84.750 ;
        RECT 112.950 84.150 113.850 84.450 ;
        RECT 118.350 84.150 119.250 84.450 ;
        RECT 112.950 83.850 114.150 84.150 ;
        RECT 118.050 83.850 119.250 84.150 ;
        RECT 32.780 82.580 37.280 83.780 ;
        RECT 112.950 83.550 114.750 83.850 ;
        RECT 117.450 83.550 119.250 83.850 ;
        RECT 112.950 83.250 115.350 83.550 ;
        RECT 116.850 83.250 118.950 83.550 ;
        RECT 111.850 82.820 112.960 83.050 ;
        RECT 114.750 82.950 115.950 83.250 ;
        RECT 116.250 82.950 117.450 83.250 ;
        RECT 32.780 82.280 33.680 82.580 ;
        RECT 32.780 81.980 33.380 82.280 ;
        RECT 33.080 81.680 33.380 81.980 ;
        RECT 34.580 81.680 35.480 82.580 ;
        RECT 36.380 82.280 37.280 82.580 ;
        RECT 36.680 81.980 37.280 82.280 ;
        RECT 110.660 82.320 112.960 82.820 ;
        RECT 115.350 82.350 116.850 82.950 ;
        RECT 119.070 82.820 120.130 83.050 ;
        RECT 120.420 82.820 120.920 95.290 ;
        RECT 121.290 94.970 122.400 95.290 ;
        RECT 124.790 95.270 126.290 95.870 ;
        RECT 128.510 95.790 130.020 95.970 ;
        RECT 128.510 95.290 130.110 95.790 ;
        RECT 124.190 94.970 125.390 95.270 ;
        RECT 125.690 94.970 126.890 95.270 ;
        RECT 128.510 94.970 129.570 95.290 ;
        RECT 123.590 94.670 124.790 94.970 ;
        RECT 126.290 94.670 127.490 94.970 ;
        RECT 122.690 94.370 124.490 94.670 ;
        RECT 126.590 94.370 128.390 94.670 ;
        RECT 122.390 93.770 123.890 94.370 ;
        RECT 127.190 93.770 128.690 94.370 ;
        RECT 122.690 93.470 123.590 93.770 ;
        RECT 124.490 93.470 124.790 93.770 ;
        RECT 125.090 93.470 125.390 93.770 ;
        RECT 125.690 93.470 125.990 93.770 ;
        RECT 126.290 93.470 126.590 93.770 ;
        RECT 127.490 93.470 128.390 93.770 ;
        RECT 124.490 92.870 126.590 93.470 ;
        RECT 123.890 92.570 125.090 92.870 ;
        RECT 125.990 92.570 126.890 92.870 ;
        RECT 123.890 92.270 125.390 92.570 ;
        RECT 125.690 92.270 127.490 92.570 ;
        RECT 123.590 91.970 124.190 92.270 ;
        RECT 124.790 91.970 126.290 92.270 ;
        RECT 126.890 91.970 127.490 92.270 ;
        RECT 123.590 91.670 123.890 91.970 ;
        RECT 123.290 91.370 123.890 91.670 ;
        RECT 123.290 91.070 124.190 91.370 ;
        RECT 125.090 91.070 125.990 91.970 ;
        RECT 127.190 91.670 127.490 91.970 ;
        RECT 127.190 91.370 127.790 91.670 ;
        RECT 126.890 91.070 127.790 91.370 ;
        RECT 123.290 89.870 127.790 91.070 ;
        RECT 123.590 89.270 127.490 89.870 ;
        RECT 124.190 88.970 126.890 89.270 ;
        RECT 127.960 89.240 129.070 89.740 ;
        RECT 128.620 89.130 129.070 89.240 ;
        RECT 124.190 88.670 126.590 88.970 ;
        RECT 36.680 81.680 36.980 81.980 ;
        RECT 33.080 81.380 33.680 81.680 ;
        RECT 34.280 81.380 35.780 81.680 ;
        RECT 36.380 81.380 36.980 81.680 ;
        RECT 33.380 81.080 34.880 81.380 ;
        RECT 35.180 81.080 36.980 81.380 ;
        RECT 33.380 80.780 34.580 81.080 ;
        RECT 35.480 80.780 36.380 81.080 ;
        RECT 33.980 80.180 36.080 80.780 ;
        RECT 32.180 79.880 32.480 80.180 ;
        RECT 33.980 79.880 34.280 80.180 ;
        RECT 34.580 79.880 34.880 80.180 ;
        RECT 35.180 79.880 35.480 80.180 ;
        RECT 35.780 79.880 36.080 80.180 ;
        RECT 37.580 79.880 37.880 80.180 ;
        RECT 31.880 79.580 32.780 79.880 ;
        RECT 37.280 79.580 38.180 79.880 ;
        RECT 31.880 79.280 33.080 79.580 ;
        RECT 36.980 79.280 38.180 79.580 ;
        RECT 31.880 78.980 33.680 79.280 ;
        RECT 36.380 78.980 38.180 79.280 ;
        RECT 104.210 79.390 106.610 79.690 ;
        RECT 104.210 79.090 106.910 79.390 ;
        RECT 108.530 79.130 109.090 79.300 ;
        RECT 31.880 78.680 34.280 78.980 ;
        RECT 35.780 78.680 37.880 78.980 ;
        RECT 30.280 77.730 31.890 78.480 ;
        RECT 33.680 78.380 34.880 78.680 ;
        RECT 35.180 78.380 36.380 78.680 ;
        RECT 103.610 78.490 107.510 79.090 ;
        RECT 107.700 78.690 109.090 79.130 ;
        RECT 34.280 77.780 35.780 78.380 ;
        RECT 38.000 78.250 39.060 78.480 ;
        RECT 38.000 78.230 39.560 78.250 ;
        RECT 30.780 77.480 31.890 77.730 ;
        RECT 33.680 77.480 34.880 77.780 ;
        RECT 35.180 77.480 36.380 77.780 ;
        RECT 38.000 77.730 41.870 78.230 ;
        RECT 38.000 77.480 39.060 77.730 ;
        RECT 33.080 77.180 34.280 77.480 ;
        RECT 35.780 77.180 36.980 77.480 ;
        RECT 32.180 76.880 33.980 77.180 ;
        RECT 36.080 76.880 37.880 77.180 ;
        RECT 31.880 76.280 33.380 76.880 ;
        RECT 36.680 76.280 38.180 76.880 ;
        RECT 32.180 75.980 33.080 76.280 ;
        RECT 33.980 75.980 34.280 76.280 ;
        RECT 34.580 75.980 34.880 76.280 ;
        RECT 35.180 75.980 35.480 76.280 ;
        RECT 35.780 75.980 36.080 76.280 ;
        RECT 36.980 75.980 37.880 76.280 ;
        RECT 33.980 75.380 36.080 75.980 ;
        RECT 33.380 75.080 34.580 75.380 ;
        RECT 35.480 75.080 36.380 75.380 ;
        RECT 33.380 74.780 34.880 75.080 ;
        RECT 35.180 74.780 36.980 75.080 ;
        RECT 33.080 74.480 33.680 74.780 ;
        RECT 34.280 74.480 35.780 74.780 ;
        RECT 36.380 74.480 36.980 74.780 ;
        RECT 33.080 74.180 33.380 74.480 ;
        RECT 32.780 73.880 33.380 74.180 ;
        RECT 32.780 73.580 33.680 73.880 ;
        RECT 34.580 73.580 35.480 74.480 ;
        RECT 36.680 74.180 36.980 74.480 ;
        RECT 36.680 73.880 37.280 74.180 ;
        RECT 36.380 73.580 37.280 73.880 ;
        RECT 32.780 72.380 37.280 73.580 ;
        RECT 33.080 71.780 36.980 72.380 ;
        RECT 33.680 71.480 36.380 71.780 ;
        RECT 37.450 71.750 38.560 72.250 ;
        RECT 38.110 71.640 38.560 71.750 ;
        RECT 33.680 71.180 36.080 71.480 ;
        RECT 41.370 68.580 41.870 77.730 ;
        RECT 103.310 77.290 107.810 78.490 ;
        RECT 103.310 76.990 104.210 77.290 ;
        RECT 103.310 76.690 103.910 76.990 ;
        RECT 103.610 76.390 103.910 76.690 ;
        RECT 105.110 76.390 106.010 77.290 ;
        RECT 106.910 76.990 107.810 77.290 ;
        RECT 107.210 76.690 107.810 76.990 ;
        RECT 107.210 76.390 107.510 76.690 ;
        RECT 103.610 76.090 104.210 76.390 ;
        RECT 104.810 76.090 106.310 76.390 ;
        RECT 106.910 76.090 107.510 76.390 ;
        RECT 103.910 75.790 105.410 76.090 ;
        RECT 105.710 75.790 107.510 76.090 ;
        RECT 103.910 75.490 105.110 75.790 ;
        RECT 106.010 75.490 106.910 75.790 ;
        RECT 45.790 75.010 48.190 75.310 ;
        RECT 45.790 74.710 48.490 75.010 ;
        RECT 50.110 74.750 50.670 74.920 ;
        RECT 104.510 74.890 106.610 75.490 ;
        RECT 45.190 74.110 49.090 74.710 ;
        RECT 49.280 74.310 50.670 74.750 ;
        RECT 102.710 74.590 103.010 74.890 ;
        RECT 104.510 74.590 104.810 74.890 ;
        RECT 105.110 74.590 105.410 74.890 ;
        RECT 105.710 74.590 106.010 74.890 ;
        RECT 106.310 74.590 106.610 74.890 ;
        RECT 108.110 74.590 108.410 74.890 ;
        RECT 102.410 74.290 103.310 74.590 ;
        RECT 107.810 74.290 108.710 74.590 ;
        RECT 44.890 72.910 49.390 74.110 ;
        RECT 102.410 73.990 103.610 74.290 ;
        RECT 107.510 73.990 108.710 74.290 ;
        RECT 102.410 73.690 104.210 73.990 ;
        RECT 106.910 73.690 108.710 73.990 ;
        RECT 102.410 73.390 104.810 73.690 ;
        RECT 106.310 73.390 108.410 73.690 ;
        RECT 101.310 72.960 102.420 73.190 ;
        RECT 104.210 73.090 105.410 73.390 ;
        RECT 105.710 73.090 106.910 73.390 ;
        RECT 100.920 72.950 102.420 72.960 ;
        RECT 44.890 72.610 45.790 72.910 ;
        RECT 44.890 72.310 45.490 72.610 ;
        RECT 45.190 72.010 45.490 72.310 ;
        RECT 46.690 72.010 47.590 72.910 ;
        RECT 48.490 72.610 49.390 72.910 ;
        RECT 48.790 72.310 49.390 72.610 ;
        RECT 98.490 72.450 102.420 72.950 ;
        RECT 104.810 72.490 106.310 73.090 ;
        RECT 108.530 72.970 109.590 73.190 ;
        RECT 110.660 72.970 111.160 82.320 ;
        RECT 111.850 82.050 112.960 82.320 ;
        RECT 114.750 82.050 115.950 82.350 ;
        RECT 116.250 82.050 117.450 82.350 ;
        RECT 119.070 82.320 120.920 82.820 ;
        RECT 119.070 82.050 120.130 82.320 ;
        RECT 120.420 82.300 120.920 82.320 ;
        RECT 114.150 81.750 115.350 82.050 ;
        RECT 116.850 81.750 118.050 82.050 ;
        RECT 113.250 81.450 115.050 81.750 ;
        RECT 117.150 81.450 118.950 81.750 ;
        RECT 112.950 80.850 114.450 81.450 ;
        RECT 117.750 80.850 119.250 81.450 ;
        RECT 113.250 80.550 114.150 80.850 ;
        RECT 115.050 80.550 115.350 80.850 ;
        RECT 115.650 80.550 115.950 80.850 ;
        RECT 116.250 80.550 116.550 80.850 ;
        RECT 116.850 80.550 117.150 80.850 ;
        RECT 118.050 80.550 118.950 80.850 ;
        RECT 115.050 79.950 117.150 80.550 ;
        RECT 114.450 79.650 115.650 79.950 ;
        RECT 116.550 79.650 117.450 79.950 ;
        RECT 114.450 79.350 115.950 79.650 ;
        RECT 116.250 79.350 118.050 79.650 ;
        RECT 114.150 79.050 114.750 79.350 ;
        RECT 115.350 79.050 116.850 79.350 ;
        RECT 117.450 79.050 118.050 79.350 ;
        RECT 114.150 78.750 114.450 79.050 ;
        RECT 113.850 78.450 114.450 78.750 ;
        RECT 113.850 78.150 114.750 78.450 ;
        RECT 115.650 78.150 116.550 79.050 ;
        RECT 117.750 78.750 118.050 79.050 ;
        RECT 117.750 78.450 118.350 78.750 ;
        RECT 117.450 78.150 118.350 78.450 ;
        RECT 113.850 76.950 118.350 78.150 ;
        RECT 114.150 76.350 118.050 76.950 ;
        RECT 114.750 76.050 117.450 76.350 ;
        RECT 118.520 76.320 119.630 76.820 ;
        RECT 119.180 76.210 119.630 76.320 ;
        RECT 114.750 75.750 117.150 76.050 ;
        RECT 48.790 72.010 49.090 72.310 ;
        RECT 45.190 71.710 45.790 72.010 ;
        RECT 46.390 71.710 47.890 72.010 ;
        RECT 48.490 71.710 49.090 72.010 ;
        RECT 45.490 71.410 46.990 71.710 ;
        RECT 47.290 71.410 49.090 71.710 ;
        RECT 90.780 71.640 93.180 71.940 ;
        RECT 45.490 71.110 46.690 71.410 ;
        RECT 47.590 71.110 48.490 71.410 ;
        RECT 90.780 71.340 93.480 71.640 ;
        RECT 95.100 71.380 95.660 71.550 ;
        RECT 46.090 70.510 48.190 71.110 ;
        RECT 90.180 70.740 94.080 71.340 ;
        RECT 94.270 70.940 95.660 71.380 ;
        RECT 44.290 70.210 44.590 70.510 ;
        RECT 46.090 70.210 46.390 70.510 ;
        RECT 46.690 70.210 46.990 70.510 ;
        RECT 47.290 70.210 47.590 70.510 ;
        RECT 47.890 70.210 48.190 70.510 ;
        RECT 49.690 70.210 49.990 70.510 ;
        RECT 43.990 69.910 44.890 70.210 ;
        RECT 49.390 69.910 50.290 70.210 ;
        RECT 43.990 69.610 45.190 69.910 ;
        RECT 49.090 69.610 50.290 69.910 ;
        RECT 43.990 69.310 45.790 69.610 ;
        RECT 48.490 69.310 50.290 69.610 ;
        RECT 60.220 69.350 62.620 69.650 ;
        RECT 89.880 69.540 94.380 70.740 ;
        RECT 43.990 69.010 46.390 69.310 ;
        RECT 47.890 69.010 49.990 69.310 ;
        RECT 60.220 69.050 62.920 69.350 ;
        RECT 64.540 69.090 65.100 69.260 ;
        RECT 42.890 68.580 44.000 68.810 ;
        RECT 45.790 68.710 46.990 69.010 ;
        RECT 47.290 68.710 48.490 69.010 ;
        RECT 41.280 68.080 44.000 68.580 ;
        RECT 46.390 68.110 47.890 68.710 ;
        RECT 50.110 68.580 51.170 68.810 ;
        RECT 50.110 68.560 51.670 68.580 ;
        RECT 42.890 67.810 44.000 68.080 ;
        RECT 45.790 67.810 46.990 68.110 ;
        RECT 47.290 67.810 48.490 68.110 ;
        RECT 50.110 68.060 54.940 68.560 ;
        RECT 59.620 68.450 63.520 69.050 ;
        RECT 63.710 68.650 65.100 69.090 ;
        RECT 89.880 69.240 90.780 69.540 ;
        RECT 89.880 68.940 90.480 69.240 ;
        RECT 90.180 68.640 90.480 68.940 ;
        RECT 91.680 68.640 92.580 69.540 ;
        RECT 93.480 69.240 94.380 69.540 ;
        RECT 93.780 68.940 94.380 69.240 ;
        RECT 93.780 68.640 94.080 68.940 ;
        RECT 50.110 67.810 51.170 68.060 ;
        RECT 45.190 67.510 46.390 67.810 ;
        RECT 47.890 67.510 49.090 67.810 ;
        RECT 44.290 67.210 46.090 67.510 ;
        RECT 48.190 67.210 49.990 67.510 ;
        RECT 43.990 66.610 45.490 67.210 ;
        RECT 48.790 66.610 50.290 67.210 ;
        RECT 44.290 66.310 45.190 66.610 ;
        RECT 46.090 66.310 46.390 66.610 ;
        RECT 46.690 66.310 46.990 66.610 ;
        RECT 47.290 66.310 47.590 66.610 ;
        RECT 47.890 66.310 48.190 66.610 ;
        RECT 49.090 66.310 49.990 66.610 ;
        RECT 46.090 65.710 48.190 66.310 ;
        RECT 45.490 65.410 46.690 65.710 ;
        RECT 47.590 65.410 48.490 65.710 ;
        RECT 45.490 65.110 46.990 65.410 ;
        RECT 47.290 65.110 49.090 65.410 ;
        RECT 45.190 64.810 45.790 65.110 ;
        RECT 46.390 64.810 47.890 65.110 ;
        RECT 48.490 64.810 49.090 65.110 ;
        RECT 45.190 64.510 45.490 64.810 ;
        RECT 44.890 64.210 45.490 64.510 ;
        RECT 44.890 63.910 45.790 64.210 ;
        RECT 46.690 63.910 47.590 64.810 ;
        RECT 48.790 64.510 49.090 64.810 ;
        RECT 48.790 64.210 49.390 64.510 ;
        RECT 48.490 63.910 49.390 64.210 ;
        RECT 44.890 62.710 49.390 63.910 ;
        RECT 54.440 62.920 54.940 68.060 ;
        RECT 59.320 67.250 63.820 68.450 ;
        RECT 75.670 68.190 78.070 68.490 ;
        RECT 90.180 68.340 90.780 68.640 ;
        RECT 91.380 68.340 92.880 68.640 ;
        RECT 93.480 68.340 94.080 68.640 ;
        RECT 75.670 67.890 78.370 68.190 ;
        RECT 79.990 67.930 80.550 68.100 ;
        RECT 75.070 67.290 78.970 67.890 ;
        RECT 79.160 67.490 80.550 67.930 ;
        RECT 90.480 68.040 91.980 68.340 ;
        RECT 92.280 68.040 94.080 68.340 ;
        RECT 90.480 67.740 91.680 68.040 ;
        RECT 92.580 67.740 93.480 68.040 ;
        RECT 59.320 66.950 60.220 67.250 ;
        RECT 59.320 66.650 59.920 66.950 ;
        RECT 59.620 66.350 59.920 66.650 ;
        RECT 61.120 66.350 62.020 67.250 ;
        RECT 62.920 66.950 63.820 67.250 ;
        RECT 63.220 66.650 63.820 66.950 ;
        RECT 63.220 66.350 63.520 66.650 ;
        RECT 59.620 66.050 60.220 66.350 ;
        RECT 60.820 66.050 62.320 66.350 ;
        RECT 62.920 66.050 63.520 66.350 ;
        RECT 59.920 65.750 61.420 66.050 ;
        RECT 61.720 65.750 63.520 66.050 ;
        RECT 74.770 66.090 79.270 67.290 ;
        RECT 91.080 67.140 93.180 67.740 ;
        RECT 89.280 66.840 89.580 67.140 ;
        RECT 91.080 66.840 91.380 67.140 ;
        RECT 91.680 66.840 91.980 67.140 ;
        RECT 92.280 66.840 92.580 67.140 ;
        RECT 92.880 66.840 93.180 67.140 ;
        RECT 94.680 66.840 94.980 67.140 ;
        RECT 74.770 65.790 75.670 66.090 ;
        RECT 59.920 65.450 61.120 65.750 ;
        RECT 62.020 65.450 62.920 65.750 ;
        RECT 74.770 65.490 75.370 65.790 ;
        RECT 60.520 64.850 62.620 65.450 ;
        RECT 75.070 65.190 75.370 65.490 ;
        RECT 76.570 65.190 77.470 66.090 ;
        RECT 78.370 65.790 79.270 66.090 ;
        RECT 78.670 65.490 79.270 65.790 ;
        RECT 88.980 66.540 89.880 66.840 ;
        RECT 94.380 66.540 95.280 66.840 ;
        RECT 88.980 66.240 90.180 66.540 ;
        RECT 94.080 66.240 95.280 66.540 ;
        RECT 88.980 65.940 90.780 66.240 ;
        RECT 93.480 65.940 95.280 66.240 ;
        RECT 88.980 65.640 91.380 65.940 ;
        RECT 92.880 65.640 94.980 65.940 ;
        RECT 78.670 65.190 78.970 65.490 ;
        RECT 87.880 65.210 88.990 65.440 ;
        RECT 90.780 65.340 91.980 65.640 ;
        RECT 92.280 65.340 93.480 65.640 ;
        RECT 75.070 64.890 75.670 65.190 ;
        RECT 76.270 64.890 77.770 65.190 ;
        RECT 78.370 64.890 78.970 65.190 ;
        RECT 58.720 64.550 59.020 64.850 ;
        RECT 60.520 64.550 60.820 64.850 ;
        RECT 61.120 64.550 61.420 64.850 ;
        RECT 61.720 64.550 62.020 64.850 ;
        RECT 62.320 64.550 62.620 64.850 ;
        RECT 64.120 64.550 64.420 64.850 ;
        RECT 75.370 64.590 76.870 64.890 ;
        RECT 77.170 64.590 78.970 64.890 ;
        RECT 84.430 64.710 88.990 65.210 ;
        RECT 91.380 64.740 92.880 65.340 ;
        RECT 95.100 65.210 96.160 65.440 ;
        RECT 98.490 65.210 98.990 72.450 ;
        RECT 101.310 72.190 102.420 72.450 ;
        RECT 104.210 72.190 105.410 72.490 ;
        RECT 105.710 72.190 106.910 72.490 ;
        RECT 108.530 72.470 111.160 72.970 ;
        RECT 108.530 72.460 110.090 72.470 ;
        RECT 108.530 72.190 109.590 72.460 ;
        RECT 103.610 71.890 104.810 72.190 ;
        RECT 106.310 71.890 107.510 72.190 ;
        RECT 102.710 71.590 104.510 71.890 ;
        RECT 106.610 71.590 108.410 71.890 ;
        RECT 102.410 70.990 103.910 71.590 ;
        RECT 107.210 70.990 108.710 71.590 ;
        RECT 102.710 70.690 103.610 70.990 ;
        RECT 104.510 70.690 104.810 70.990 ;
        RECT 105.110 70.690 105.410 70.990 ;
        RECT 105.710 70.690 106.010 70.990 ;
        RECT 106.310 70.690 106.610 70.990 ;
        RECT 107.510 70.690 108.410 70.990 ;
        RECT 104.510 70.090 106.610 70.690 ;
        RECT 103.910 69.790 105.110 70.090 ;
        RECT 106.010 69.790 106.910 70.090 ;
        RECT 103.910 69.490 105.410 69.790 ;
        RECT 105.710 69.490 107.510 69.790 ;
        RECT 103.610 69.190 104.210 69.490 ;
        RECT 104.810 69.190 106.310 69.490 ;
        RECT 106.910 69.190 107.510 69.490 ;
        RECT 103.610 68.890 103.910 69.190 ;
        RECT 103.310 68.590 103.910 68.890 ;
        RECT 103.310 68.290 104.210 68.590 ;
        RECT 105.110 68.290 106.010 69.190 ;
        RECT 107.210 68.890 107.510 69.190 ;
        RECT 107.210 68.590 107.810 68.890 ;
        RECT 106.910 68.290 107.810 68.590 ;
        RECT 103.310 67.090 107.810 68.290 ;
        RECT 103.610 66.490 107.510 67.090 ;
        RECT 104.210 66.190 106.910 66.490 ;
        RECT 107.980 66.460 109.090 66.960 ;
        RECT 108.640 66.350 109.090 66.460 ;
        RECT 104.210 65.890 106.610 66.190 ;
        RECT 58.420 64.250 59.320 64.550 ;
        RECT 63.820 64.250 64.720 64.550 ;
        RECT 75.370 64.290 76.570 64.590 ;
        RECT 77.470 64.290 78.370 64.590 ;
        RECT 58.420 63.950 59.620 64.250 ;
        RECT 63.520 63.950 64.720 64.250 ;
        RECT 58.420 63.650 60.220 63.950 ;
        RECT 62.920 63.650 64.720 63.950 ;
        RECT 75.970 63.690 78.070 64.290 ;
        RECT 58.420 63.350 60.820 63.650 ;
        RECT 62.320 63.350 64.420 63.650 ;
        RECT 74.170 63.390 74.470 63.690 ;
        RECT 75.970 63.390 76.270 63.690 ;
        RECT 76.570 63.390 76.870 63.690 ;
        RECT 77.170 63.390 77.470 63.690 ;
        RECT 77.770 63.390 78.070 63.690 ;
        RECT 79.570 63.390 79.870 63.690 ;
        RECT 57.320 62.920 58.430 63.150 ;
        RECT 60.220 63.050 61.420 63.350 ;
        RECT 61.720 63.050 62.920 63.350 ;
        RECT 45.190 62.110 49.090 62.710 ;
        RECT 45.790 61.810 48.490 62.110 ;
        RECT 49.560 62.080 50.670 62.580 ;
        RECT 54.440 62.420 58.430 62.920 ;
        RECT 60.820 62.450 62.320 63.050 ;
        RECT 64.540 62.940 65.600 63.150 ;
        RECT 73.870 63.090 74.770 63.390 ;
        RECT 79.270 63.090 80.170 63.390 ;
        RECT 57.320 62.150 58.430 62.420 ;
        RECT 60.220 62.150 61.420 62.450 ;
        RECT 61.720 62.150 62.920 62.450 ;
        RECT 64.540 62.440 69.780 62.940 ;
        RECT 64.540 62.420 66.100 62.440 ;
        RECT 64.540 62.150 65.600 62.420 ;
        RECT 50.220 61.970 50.670 62.080 ;
        RECT 59.620 61.850 60.820 62.150 ;
        RECT 62.320 61.850 63.520 62.150 ;
        RECT 45.790 61.510 48.190 61.810 ;
        RECT 58.720 61.550 60.520 61.850 ;
        RECT 62.620 61.550 64.420 61.850 ;
        RECT 69.280 61.760 69.780 62.440 ;
        RECT 73.870 62.790 75.070 63.090 ;
        RECT 78.970 62.790 80.170 63.090 ;
        RECT 73.870 62.490 75.670 62.790 ;
        RECT 78.370 62.490 80.170 62.790 ;
        RECT 73.870 62.190 76.270 62.490 ;
        RECT 77.770 62.190 79.870 62.490 ;
        RECT 72.770 61.760 73.880 61.990 ;
        RECT 75.670 61.890 76.870 62.190 ;
        RECT 77.170 61.890 78.370 62.190 ;
        RECT 58.420 60.950 59.920 61.550 ;
        RECT 63.220 60.950 64.720 61.550 ;
        RECT 69.280 61.260 73.880 61.760 ;
        RECT 76.270 61.290 77.770 61.890 ;
        RECT 79.990 61.760 81.050 61.990 ;
        RECT 79.990 61.720 81.550 61.760 ;
        RECT 84.430 61.720 84.930 64.710 ;
        RECT 87.880 64.440 88.990 64.710 ;
        RECT 90.780 64.440 91.980 64.740 ;
        RECT 92.280 64.440 93.480 64.740 ;
        RECT 95.100 64.710 98.990 65.210 ;
        RECT 95.100 64.440 96.160 64.710 ;
        RECT 90.180 64.140 91.380 64.440 ;
        RECT 92.880 64.140 94.080 64.440 ;
        RECT 89.280 63.840 91.080 64.140 ;
        RECT 93.180 63.840 94.980 64.140 ;
        RECT 88.980 63.240 90.480 63.840 ;
        RECT 93.780 63.240 95.280 63.840 ;
        RECT 89.280 62.940 90.180 63.240 ;
        RECT 91.080 62.940 91.380 63.240 ;
        RECT 91.680 62.940 91.980 63.240 ;
        RECT 92.280 62.940 92.580 63.240 ;
        RECT 92.880 62.940 93.180 63.240 ;
        RECT 94.080 62.940 94.980 63.240 ;
        RECT 91.080 62.340 93.180 62.940 ;
        RECT 90.480 62.040 91.680 62.340 ;
        RECT 92.580 62.040 93.480 62.340 ;
        RECT 90.480 61.740 91.980 62.040 ;
        RECT 92.280 61.740 94.080 62.040 ;
        RECT 72.770 60.990 73.880 61.260 ;
        RECT 75.670 60.990 76.870 61.290 ;
        RECT 77.170 60.990 78.370 61.290 ;
        RECT 79.990 61.220 84.930 61.720 ;
        RECT 90.180 61.440 90.780 61.740 ;
        RECT 91.380 61.440 92.880 61.740 ;
        RECT 93.480 61.440 94.080 61.740 ;
        RECT 79.990 60.990 81.050 61.220 ;
        RECT 90.180 61.140 90.480 61.440 ;
        RECT 58.720 60.650 59.620 60.950 ;
        RECT 60.520 60.650 60.820 60.950 ;
        RECT 61.120 60.650 61.420 60.950 ;
        RECT 61.720 60.650 62.020 60.950 ;
        RECT 62.320 60.650 62.620 60.950 ;
        RECT 63.520 60.650 64.420 60.950 ;
        RECT 75.070 60.690 76.270 60.990 ;
        RECT 77.770 60.690 78.970 60.990 ;
        RECT 89.880 60.840 90.480 61.140 ;
        RECT 60.520 60.050 62.620 60.650 ;
        RECT 74.170 60.390 75.970 60.690 ;
        RECT 78.070 60.390 79.870 60.690 ;
        RECT 89.880 60.540 90.780 60.840 ;
        RECT 91.680 60.540 92.580 61.440 ;
        RECT 93.780 61.140 94.080 61.440 ;
        RECT 93.780 60.840 94.380 61.140 ;
        RECT 93.480 60.540 94.380 60.840 ;
        RECT 59.920 59.750 61.120 60.050 ;
        RECT 62.020 59.750 62.920 60.050 ;
        RECT 73.870 59.790 75.370 60.390 ;
        RECT 78.670 59.790 80.170 60.390 ;
        RECT 59.920 59.450 61.420 59.750 ;
        RECT 61.720 59.450 63.520 59.750 ;
        RECT 74.170 59.490 75.070 59.790 ;
        RECT 75.970 59.490 76.270 59.790 ;
        RECT 76.570 59.490 76.870 59.790 ;
        RECT 77.170 59.490 77.470 59.790 ;
        RECT 77.770 59.490 78.070 59.790 ;
        RECT 78.970 59.490 79.870 59.790 ;
        RECT 59.620 59.150 60.220 59.450 ;
        RECT 60.820 59.150 62.320 59.450 ;
        RECT 62.920 59.150 63.520 59.450 ;
        RECT 59.620 58.850 59.920 59.150 ;
        RECT 59.320 58.550 59.920 58.850 ;
        RECT 59.320 58.250 60.220 58.550 ;
        RECT 61.120 58.250 62.020 59.150 ;
        RECT 63.220 58.850 63.520 59.150 ;
        RECT 75.970 58.890 78.070 59.490 ;
        RECT 89.880 59.340 94.380 60.540 ;
        RECT 63.220 58.550 63.820 58.850 ;
        RECT 62.920 58.250 63.820 58.550 ;
        RECT 75.370 58.590 76.570 58.890 ;
        RECT 77.470 58.590 78.370 58.890 ;
        RECT 90.180 58.740 94.080 59.340 ;
        RECT 75.370 58.290 76.870 58.590 ;
        RECT 77.170 58.290 78.970 58.590 ;
        RECT 59.320 57.050 63.820 58.250 ;
        RECT 75.070 57.990 75.670 58.290 ;
        RECT 76.270 57.990 77.770 58.290 ;
        RECT 78.370 57.990 78.970 58.290 ;
        RECT 90.780 58.440 93.480 58.740 ;
        RECT 94.550 58.710 95.660 59.210 ;
        RECT 95.210 58.600 95.660 58.710 ;
        RECT 90.780 58.140 93.180 58.440 ;
        RECT 75.070 57.690 75.370 57.990 ;
        RECT 74.770 57.390 75.370 57.690 ;
        RECT 74.770 57.090 75.670 57.390 ;
        RECT 76.570 57.090 77.470 57.990 ;
        RECT 78.670 57.690 78.970 57.990 ;
        RECT 78.670 57.390 79.270 57.690 ;
        RECT 78.370 57.090 79.270 57.390 ;
        RECT 59.620 56.450 63.520 57.050 ;
        RECT 60.220 56.150 62.920 56.450 ;
        RECT 63.990 56.420 65.100 56.920 ;
        RECT 64.650 56.310 65.100 56.420 ;
        RECT 60.220 55.850 62.620 56.150 ;
        RECT 74.770 55.890 79.270 57.090 ;
        RECT 75.070 55.290 78.970 55.890 ;
        RECT 75.670 54.990 78.370 55.290 ;
        RECT 79.440 55.260 80.550 55.760 ;
        RECT 80.100 55.150 80.550 55.260 ;
        RECT 75.670 54.690 78.070 54.990 ;
      LAYER met2 ;
        RECT 70.220 223.640 70.540 224.140 ;
        RECT 72.980 223.640 73.300 224.140 ;
        RECT 70.230 222.770 70.490 223.640 ;
        RECT 48.690 222.510 70.490 222.770 ;
        RECT 48.690 219.110 48.950 222.510 ;
        RECT 73.000 222.250 73.260 223.640 ;
        RECT 58.400 221.990 73.260 222.250 ;
        RECT 48.680 218.750 48.990 219.110 ;
        RECT 58.400 219.070 58.660 221.990 ;
        RECT 75.740 221.830 76.060 224.140 ;
        RECT 68.040 221.570 76.060 221.830 ;
        RECT 68.040 219.170 68.300 221.570 ;
        RECT 76.130 220.815 76.610 221.395 ;
        RECT 74.660 219.355 75.120 220.010 ;
        RECT 45.770 218.030 46.460 218.730 ;
        RECT 58.350 218.710 58.660 219.070 ;
        RECT 67.990 218.810 68.300 219.170 ;
        RECT 44.460 215.395 45.010 215.775 ;
        RECT 36.560 215.130 37.060 215.235 ;
        RECT 51.570 215.130 52.130 216.740 ;
        RECT 36.560 214.680 39.010 215.130 ;
        RECT 36.560 214.635 37.060 214.680 ;
        RECT 43.040 214.450 43.640 214.750 ;
        RECT 45.740 214.450 46.640 214.750 ;
        RECT 50.740 214.570 52.130 215.130 ;
        RECT 39.140 213.550 40.940 213.850 ;
        RECT 42.740 213.550 43.940 214.450 ;
        RECT 45.440 214.150 46.940 214.450 ;
        RECT 45.440 213.850 46.640 214.150 ;
        RECT 45.440 213.550 46.340 213.850 ;
        RECT 48.740 213.550 50.540 213.850 ;
        RECT 38.540 213.250 41.840 213.550 ;
        RECT 43.040 213.250 44.240 213.550 ;
        RECT 38.540 212.950 40.640 213.250 ;
        RECT 41.240 212.950 41.840 213.250 ;
        RECT 43.640 212.950 44.240 213.250 ;
        RECT 45.440 212.950 46.040 213.550 ;
        RECT 47.840 213.250 51.140 213.550 ;
        RECT 47.840 212.950 48.440 213.250 ;
        RECT 49.040 212.950 51.140 213.250 ;
        RECT 38.240 212.650 40.340 212.950 ;
        RECT 37.940 212.050 40.340 212.650 ;
        RECT 41.540 212.650 42.140 212.950 ;
        RECT 43.640 212.650 44.540 212.950 ;
        RECT 41.540 212.350 43.040 212.650 ;
        RECT 43.940 212.350 44.540 212.650 ;
        RECT 45.140 212.350 45.740 212.950 ;
        RECT 47.540 212.650 48.140 212.950 ;
        RECT 46.640 212.350 48.140 212.650 ;
        RECT 49.340 212.650 51.440 212.950 ;
        RECT 41.240 212.050 42.740 212.350 ;
        RECT 37.940 211.750 41.840 212.050 ;
        RECT 42.140 211.750 43.040 212.050 ;
        RECT 44.240 211.750 45.440 212.350 ;
        RECT 46.940 212.050 48.440 212.350 ;
        RECT 49.340 212.050 51.740 212.650 ;
        RECT 46.640 211.750 47.540 212.050 ;
        RECT 47.840 211.750 51.740 212.050 ;
        RECT 37.940 211.450 41.540 211.750 ;
        RECT 42.140 211.450 42.740 211.750 ;
        RECT 44.540 211.450 45.140 211.750 ;
        RECT 46.940 211.450 47.540 211.750 ;
        RECT 48.140 211.450 51.740 211.750 ;
        RECT 37.940 211.150 41.840 211.450 ;
        RECT 42.140 211.150 43.040 211.450 ;
        RECT 37.940 210.250 40.340 211.150 ;
        RECT 41.240 210.850 42.740 211.150 ;
        RECT 44.240 210.850 45.440 211.450 ;
        RECT 46.640 211.150 47.540 211.450 ;
        RECT 47.840 211.150 51.740 211.450 ;
        RECT 46.940 210.850 48.440 211.150 ;
        RECT 41.540 210.550 43.040 210.850 ;
        RECT 43.940 210.550 44.540 210.850 ;
        RECT 41.540 210.250 42.140 210.550 ;
        RECT 38.540 209.950 40.640 210.250 ;
        RECT 41.240 209.950 42.140 210.250 ;
        RECT 43.640 210.250 44.540 210.550 ;
        RECT 45.140 210.250 45.740 210.850 ;
        RECT 46.640 210.550 48.140 210.850 ;
        RECT 47.540 210.250 48.140 210.550 ;
        RECT 49.340 210.250 51.740 211.150 ;
        RECT 43.640 209.950 44.240 210.250 ;
        RECT 38.540 209.650 41.540 209.950 ;
        RECT 43.040 209.650 44.240 209.950 ;
        RECT 45.440 209.650 46.040 210.250 ;
        RECT 47.540 209.950 48.440 210.250 ;
        RECT 49.040 209.950 51.140 210.250 ;
        RECT 48.140 209.650 51.140 209.950 ;
        RECT 39.140 209.350 40.940 209.650 ;
        RECT 42.740 208.750 43.940 209.650 ;
        RECT 45.440 209.350 46.340 209.650 ;
        RECT 48.740 209.350 50.540 209.650 ;
        RECT 45.440 209.050 46.640 209.350 ;
        RECT 45.440 208.750 46.940 209.050 ;
        RECT 43.040 208.450 43.640 208.750 ;
        RECT 45.440 208.450 46.640 208.750 ;
        RECT 73.445 178.960 75.440 178.970 ;
        RECT 72.645 178.945 76.235 178.960 ;
        RECT 71.850 178.920 77.030 178.945 ;
        RECT 71.055 178.885 77.825 178.920 ;
        RECT 70.260 178.840 78.620 178.885 ;
        RECT 69.465 178.785 79.415 178.840 ;
        RECT 68.670 178.725 80.210 178.785 ;
        RECT 67.875 178.650 81.005 178.725 ;
        RECT 67.085 178.565 81.795 178.650 ;
        RECT 66.290 178.470 82.590 178.565 ;
        RECT 65.500 178.365 83.380 178.470 ;
        RECT 64.710 178.250 84.170 178.365 ;
        RECT 63.925 178.125 84.955 178.250 ;
        RECT 63.140 177.990 85.740 178.125 ;
        RECT 62.355 177.845 86.525 177.990 ;
        RECT 61.570 177.690 87.310 177.845 ;
        RECT 60.790 177.525 88.090 177.690 ;
        RECT 60.010 177.355 88.870 177.525 ;
        RECT 59.235 177.170 89.645 177.355 ;
        RECT 58.460 176.975 90.420 177.170 ;
        RECT 57.685 176.960 91.195 176.975 ;
        RECT 57.685 176.945 73.850 176.960 ;
        RECT 75.030 176.945 91.195 176.960 ;
        RECT 57.685 176.920 73.055 176.945 ;
        RECT 75.825 176.920 91.195 176.945 ;
        RECT 57.685 176.885 72.260 176.920 ;
        RECT 76.090 176.885 91.195 176.920 ;
        RECT 57.685 176.840 71.465 176.885 ;
        RECT 57.685 176.785 70.670 176.840 ;
        RECT 57.685 176.775 69.875 176.785 ;
        RECT 56.915 176.725 69.875 176.775 ;
        RECT 56.915 176.650 69.085 176.725 ;
        RECT 56.915 176.565 68.290 176.650 ;
        RECT 76.090 176.645 76.775 176.885 ;
        RECT 77.415 176.840 91.195 176.885 ;
        RECT 78.210 176.785 91.195 176.840 ;
        RECT 79.005 176.775 91.195 176.785 ;
        RECT 79.005 176.725 91.965 176.775 ;
        RECT 79.795 176.650 91.965 176.725 ;
        RECT 56.915 176.560 67.500 176.565 ;
        RECT 56.150 176.470 67.500 176.560 ;
        RECT 56.150 176.365 66.710 176.470 ;
        RECT 56.150 176.340 65.925 176.365 ;
        RECT 55.385 176.250 65.925 176.340 ;
        RECT 55.385 176.125 65.140 176.250 ;
        RECT 55.385 176.110 64.355 176.125 ;
        RECT 54.620 175.990 64.355 176.110 ;
        RECT 54.620 175.865 63.570 175.990 ;
        RECT 53.865 175.845 63.570 175.865 ;
        RECT 53.865 175.690 62.790 175.845 ;
        RECT 53.865 175.615 62.010 175.690 ;
        RECT 53.110 175.525 62.010 175.615 ;
        RECT 53.110 175.355 61.235 175.525 ;
        RECT 52.355 175.170 60.460 175.355 ;
        RECT 52.355 175.085 59.685 175.170 ;
        RECT 51.605 174.975 59.685 175.085 ;
        RECT 51.605 174.805 58.915 174.975 ;
        RECT 50.860 174.775 58.915 174.805 ;
        RECT 50.860 174.560 58.150 174.775 ;
        RECT 50.860 174.520 57.385 174.560 ;
        RECT 50.120 174.340 57.385 174.520 ;
        RECT 50.120 174.220 56.620 174.340 ;
        RECT 49.380 174.110 56.620 174.220 ;
        RECT 49.380 173.915 55.865 174.110 ;
        RECT 48.645 173.865 55.865 173.915 ;
        RECT 48.645 173.615 55.110 173.865 ;
        RECT 48.645 173.595 54.355 173.615 ;
        RECT 47.915 173.355 54.355 173.595 ;
        RECT 47.915 173.270 53.605 173.355 ;
        RECT 47.190 173.085 53.605 173.270 ;
        RECT 47.190 172.935 52.860 173.085 ;
        RECT 46.465 172.805 52.860 172.935 ;
        RECT 46.465 172.595 52.120 172.805 ;
        RECT 45.745 172.520 52.120 172.595 ;
        RECT 45.745 172.240 51.380 172.520 ;
        RECT 60.640 172.300 61.090 175.355 ;
        RECT 76.090 173.460 76.540 176.645 ;
        RECT 80.590 176.565 91.965 176.650 ;
        RECT 81.380 176.560 91.965 176.565 ;
        RECT 81.380 176.470 92.730 176.560 ;
        RECT 82.170 176.365 92.730 176.470 ;
        RECT 82.955 176.340 92.730 176.365 ;
        RECT 82.955 176.250 93.495 176.340 ;
        RECT 83.740 176.125 93.495 176.250 ;
        RECT 84.525 176.110 93.495 176.125 ;
        RECT 84.525 175.990 94.260 176.110 ;
        RECT 85.310 175.865 94.260 175.990 ;
        RECT 85.310 175.845 95.015 175.865 ;
        RECT 86.090 175.690 95.015 175.845 ;
        RECT 86.870 175.615 95.015 175.690 ;
        RECT 86.870 175.525 95.770 175.615 ;
        RECT 87.645 175.355 95.770 175.525 ;
        RECT 88.420 175.170 96.525 175.355 ;
        RECT 89.195 175.085 96.525 175.170 ;
        RECT 89.195 174.975 97.275 175.085 ;
        RECT 89.965 174.805 97.275 174.975 ;
        RECT 89.965 174.775 98.020 174.805 ;
        RECT 90.730 174.560 98.020 174.775 ;
        RECT 78.570 174.230 80.970 174.530 ;
        RECT 78.270 173.930 80.970 174.230 ;
        RECT 91.200 174.520 98.020 174.560 ;
        RECT 91.200 174.340 98.760 174.520 ;
        RECT 63.120 173.070 65.520 173.370 ;
        RECT 77.670 173.330 81.570 173.930 ;
        RECT 62.820 172.770 65.520 173.070 ;
        RECT 45.035 172.220 51.380 172.240 ;
        RECT 45.035 171.915 50.645 172.220 ;
        RECT 62.220 172.170 66.120 172.770 ;
        RECT 45.035 171.880 49.915 171.915 ;
        RECT 44.325 171.595 49.915 171.880 ;
        RECT 44.325 171.510 49.190 171.595 ;
        RECT 43.620 171.270 49.190 171.510 ;
        RECT 43.620 171.130 48.465 171.270 ;
        RECT 42.920 170.935 48.465 171.130 ;
        RECT 61.920 170.970 66.420 172.170 ;
        RECT 77.370 172.130 81.870 173.330 ;
        RECT 77.370 171.830 78.270 172.130 ;
        RECT 77.370 171.530 77.970 171.830 ;
        RECT 42.920 170.740 47.745 170.935 ;
        RECT 42.225 170.595 47.745 170.740 ;
        RECT 61.920 170.670 62.820 170.970 ;
        RECT 42.225 170.345 47.035 170.595 ;
        RECT 61.920 170.370 62.520 170.670 ;
        RECT 41.535 170.240 47.035 170.345 ;
        RECT 41.535 169.940 46.670 170.240 ;
        RECT 40.850 169.880 46.670 169.940 ;
        RECT 40.850 169.525 45.620 169.880 ;
        RECT 40.165 169.510 45.620 169.525 ;
        RECT 40.165 169.130 44.920 169.510 ;
        RECT 40.165 169.105 44.225 169.130 ;
        RECT 39.495 168.740 44.225 169.105 ;
        RECT 39.495 168.675 43.535 168.740 ;
        RECT 38.825 168.345 43.535 168.675 ;
        RECT 38.825 168.235 42.850 168.345 ;
        RECT 38.160 167.940 42.850 168.235 ;
        RECT 38.160 167.785 42.165 167.940 ;
        RECT 37.500 167.525 42.165 167.785 ;
        RECT 37.500 167.330 41.495 167.525 ;
        RECT 36.845 167.105 41.495 167.330 ;
        RECT 36.845 166.865 40.825 167.105 ;
        RECT 36.200 166.675 40.825 166.865 ;
        RECT 36.200 166.395 40.160 166.675 ;
        RECT 46.220 166.640 46.670 169.880 ;
        RECT 62.220 170.070 62.520 170.370 ;
        RECT 63.720 170.070 64.620 170.970 ;
        RECT 65.520 170.670 66.420 170.970 ;
        RECT 65.820 170.370 66.420 170.670 ;
        RECT 77.670 171.230 77.970 171.530 ;
        RECT 79.170 171.230 80.070 172.130 ;
        RECT 80.970 171.830 81.870 172.130 ;
        RECT 81.270 171.530 81.870 171.830 ;
        RECT 81.270 171.230 81.570 171.530 ;
        RECT 77.670 170.930 78.270 171.230 ;
        RECT 78.870 170.930 80.370 171.230 ;
        RECT 80.970 170.930 81.570 171.230 ;
        RECT 77.670 170.630 79.470 170.930 ;
        RECT 79.770 170.630 81.270 170.930 ;
        RECT 65.820 170.070 66.120 170.370 ;
        RECT 78.270 170.330 79.170 170.630 ;
        RECT 80.070 170.330 81.270 170.630 ;
        RECT 62.220 169.770 62.820 170.070 ;
        RECT 63.420 169.770 64.920 170.070 ;
        RECT 65.520 169.770 66.120 170.070 ;
        RECT 62.220 169.470 64.020 169.770 ;
        RECT 64.320 169.470 65.820 169.770 ;
        RECT 78.570 169.730 80.670 170.330 ;
        RECT 91.200 170.010 91.650 174.340 ;
        RECT 92.260 174.220 98.760 174.340 ;
        RECT 92.260 174.110 99.500 174.220 ;
        RECT 93.015 173.915 99.500 174.110 ;
        RECT 93.015 173.865 100.235 173.915 ;
        RECT 93.770 173.615 100.235 173.865 ;
        RECT 94.525 173.595 100.235 173.615 ;
        RECT 94.525 173.355 100.965 173.595 ;
        RECT 95.275 173.270 100.965 173.355 ;
        RECT 95.275 173.085 101.690 173.270 ;
        RECT 96.020 172.935 101.690 173.085 ;
        RECT 96.020 172.805 102.415 172.935 ;
        RECT 96.760 172.595 102.415 172.805 ;
        RECT 96.760 172.520 103.135 172.595 ;
        RECT 97.500 172.240 103.135 172.520 ;
        RECT 97.500 172.220 103.845 172.240 ;
        RECT 98.235 171.915 103.845 172.220 ;
        RECT 98.965 171.880 103.845 171.915 ;
        RECT 98.965 171.595 104.555 171.880 ;
        RECT 99.690 171.510 104.555 171.595 ;
        RECT 99.690 171.270 105.260 171.510 ;
        RECT 100.415 171.130 105.260 171.270 ;
        RECT 93.680 170.780 96.080 171.080 ;
        RECT 100.415 170.935 105.960 171.130 ;
        RECT 93.380 170.480 96.080 170.780 ;
        RECT 101.135 170.740 105.960 170.935 ;
        RECT 101.135 170.595 106.655 170.740 ;
        RECT 92.780 169.880 96.680 170.480 ;
        RECT 101.845 170.345 106.655 170.595 ;
        RECT 101.845 170.240 107.345 170.345 ;
        RECT 102.555 169.940 107.345 170.240 ;
        RECT 102.555 169.880 108.030 169.940 ;
        RECT 62.820 169.170 63.720 169.470 ;
        RECT 64.620 169.170 65.820 169.470 ;
        RECT 76.770 169.430 77.670 169.730 ;
        RECT 78.570 169.430 78.870 169.730 ;
        RECT 79.170 169.430 79.470 169.730 ;
        RECT 79.770 169.430 80.070 169.730 ;
        RECT 80.370 169.430 80.670 169.730 ;
        RECT 81.570 169.430 82.470 169.730 ;
        RECT 63.120 168.570 65.220 169.170 ;
        RECT 76.470 168.830 77.970 169.430 ;
        RECT 81.270 168.830 82.770 169.430 ;
        RECT 61.320 168.270 62.220 168.570 ;
        RECT 63.120 168.270 63.420 168.570 ;
        RECT 63.720 168.270 64.020 168.570 ;
        RECT 64.320 168.270 64.620 168.570 ;
        RECT 64.920 168.270 65.220 168.570 ;
        RECT 66.120 168.270 67.020 168.570 ;
        RECT 76.770 168.530 78.570 168.830 ;
        RECT 80.670 168.530 82.470 168.830 ;
        RECT 92.480 168.680 96.980 169.880 ;
        RECT 103.260 169.525 108.030 169.880 ;
        RECT 103.260 169.510 108.715 169.525 ;
        RECT 103.960 169.130 108.715 169.510 ;
        RECT 48.700 167.410 51.100 167.710 ;
        RECT 61.020 167.670 62.520 168.270 ;
        RECT 65.820 167.670 67.320 168.270 ;
        RECT 77.670 168.230 78.870 168.530 ;
        RECT 80.370 168.230 81.570 168.530 ;
        RECT 92.480 168.380 93.380 168.680 ;
        RECT 78.270 167.930 79.470 168.230 ;
        RECT 79.770 167.930 80.970 168.230 ;
        RECT 92.480 168.080 93.080 168.380 ;
        RECT 48.400 167.110 51.100 167.410 ;
        RECT 61.320 167.370 63.120 167.670 ;
        RECT 65.220 167.370 67.020 167.670 ;
        RECT 47.800 166.510 51.700 167.110 ;
        RECT 62.220 167.070 63.420 167.370 ;
        RECT 64.920 167.070 66.120 167.370 ;
        RECT 78.870 167.330 80.370 167.930 ;
        RECT 92.780 167.780 93.080 168.080 ;
        RECT 94.280 167.780 95.180 168.680 ;
        RECT 96.080 168.380 96.980 168.680 ;
        RECT 96.380 168.080 96.980 168.380 ;
        RECT 104.630 169.105 108.715 169.130 ;
        RECT 104.630 168.740 109.385 169.105 ;
        RECT 96.380 167.780 96.680 168.080 ;
        RECT 92.780 167.480 93.380 167.780 ;
        RECT 93.980 167.480 95.480 167.780 ;
        RECT 96.080 167.480 96.680 167.780 ;
        RECT 62.820 166.770 64.020 167.070 ;
        RECT 64.320 166.770 65.520 167.070 ;
        RECT 78.270 167.030 79.470 167.330 ;
        RECT 79.770 167.030 80.970 167.330 ;
        RECT 92.780 167.180 94.580 167.480 ;
        RECT 94.880 167.180 96.380 167.480 ;
        RECT 35.560 166.235 40.160 166.395 ;
        RECT 35.560 165.915 39.500 166.235 ;
        RECT 34.925 165.785 39.500 165.915 ;
        RECT 34.925 165.425 38.845 165.785 ;
        RECT 34.295 165.330 38.845 165.425 ;
        RECT 34.295 164.930 38.200 165.330 ;
        RECT 33.670 164.865 38.200 164.930 ;
        RECT 47.500 165.310 52.000 166.510 ;
        RECT 63.420 166.170 64.920 166.770 ;
        RECT 76.770 166.730 78.870 167.030 ;
        RECT 80.370 166.730 82.770 167.030 ;
        RECT 93.380 166.880 94.280 167.180 ;
        RECT 95.180 166.880 96.380 167.180 ;
        RECT 76.470 166.430 78.270 166.730 ;
        RECT 80.970 166.430 82.770 166.730 ;
        RECT 62.820 165.870 64.020 166.170 ;
        RECT 64.320 165.870 65.520 166.170 ;
        RECT 76.470 166.130 77.670 166.430 ;
        RECT 81.570 166.130 82.770 166.430 ;
        RECT 93.680 166.280 95.780 166.880 ;
        RECT 61.320 165.570 63.420 165.870 ;
        RECT 64.920 165.570 67.320 165.870 ;
        RECT 76.470 165.830 77.370 166.130 ;
        RECT 81.870 165.830 82.770 166.130 ;
        RECT 91.880 165.980 92.780 166.280 ;
        RECT 93.680 165.980 93.980 166.280 ;
        RECT 94.280 165.980 94.580 166.280 ;
        RECT 94.880 165.980 95.180 166.280 ;
        RECT 95.480 165.980 95.780 166.280 ;
        RECT 96.680 165.980 97.580 166.280 ;
        RECT 47.500 165.010 48.400 165.310 ;
        RECT 33.670 164.425 37.560 164.865 ;
        RECT 47.500 164.710 48.100 165.010 ;
        RECT 33.055 164.395 37.560 164.425 ;
        RECT 47.800 164.410 48.100 164.710 ;
        RECT 49.300 164.410 50.200 165.310 ;
        RECT 51.100 165.010 52.000 165.310 ;
        RECT 51.400 164.710 52.000 165.010 ;
        RECT 61.020 165.270 62.820 165.570 ;
        RECT 65.520 165.270 67.320 165.570 ;
        RECT 76.770 165.530 77.070 165.830 ;
        RECT 78.570 165.530 78.870 165.830 ;
        RECT 79.170 165.530 79.470 165.830 ;
        RECT 79.770 165.530 80.070 165.830 ;
        RECT 80.370 165.530 80.670 165.830 ;
        RECT 82.170 165.530 82.470 165.830 ;
        RECT 61.020 164.970 62.220 165.270 ;
        RECT 66.120 164.970 67.320 165.270 ;
        RECT 51.400 164.410 51.700 164.710 ;
        RECT 61.020 164.670 61.920 164.970 ;
        RECT 66.420 164.670 67.320 164.970 ;
        RECT 78.570 164.930 80.670 165.530 ;
        RECT 91.580 165.380 93.080 165.980 ;
        RECT 96.380 165.380 97.880 165.980 ;
        RECT 91.880 165.080 93.680 165.380 ;
        RECT 95.780 165.080 97.580 165.380 ;
        RECT 33.055 163.915 36.925 164.395 ;
        RECT 47.800 164.110 48.400 164.410 ;
        RECT 49.000 164.110 50.500 164.410 ;
        RECT 51.100 164.110 51.700 164.410 ;
        RECT 61.320 164.370 61.620 164.670 ;
        RECT 63.120 164.370 63.420 164.670 ;
        RECT 63.720 164.370 64.020 164.670 ;
        RECT 64.320 164.370 64.620 164.670 ;
        RECT 64.920 164.370 65.220 164.670 ;
        RECT 66.720 164.370 67.020 164.670 ;
        RECT 78.270 164.630 79.170 164.930 ;
        RECT 80.070 164.630 81.270 164.930 ;
        RECT 92.780 164.780 93.980 165.080 ;
        RECT 95.480 164.780 96.680 165.080 ;
        RECT 32.445 163.425 36.295 163.915 ;
        RECT 47.800 163.810 49.600 164.110 ;
        RECT 49.900 163.810 51.400 164.110 ;
        RECT 48.400 163.510 49.300 163.810 ;
        RECT 50.200 163.510 51.400 163.810 ;
        RECT 63.120 163.770 65.220 164.370 ;
        RECT 77.670 164.330 79.470 164.630 ;
        RECT 79.770 164.330 81.270 164.630 ;
        RECT 93.380 164.480 94.580 164.780 ;
        RECT 94.880 164.480 96.080 164.780 ;
        RECT 77.670 164.030 78.270 164.330 ;
        RECT 78.870 164.030 80.370 164.330 ;
        RECT 80.970 164.030 81.570 164.330 ;
        RECT 32.445 163.395 35.670 163.425 ;
        RECT 31.840 162.930 35.670 163.395 ;
        RECT 31.840 162.870 35.055 162.930 ;
        RECT 48.700 162.910 50.800 163.510 ;
        RECT 62.820 163.470 63.720 163.770 ;
        RECT 64.620 163.470 65.820 163.770 ;
        RECT 77.670 163.730 77.970 164.030 ;
        RECT 62.220 163.170 64.020 163.470 ;
        RECT 64.320 163.170 65.820 163.470 ;
        RECT 77.370 163.430 77.970 163.730 ;
        RECT 31.245 162.425 35.055 162.870 ;
        RECT 46.900 162.610 47.800 162.910 ;
        RECT 48.700 162.610 49.000 162.910 ;
        RECT 49.300 162.610 49.600 162.910 ;
        RECT 49.900 162.610 50.200 162.910 ;
        RECT 50.500 162.610 50.800 162.910 ;
        RECT 51.700 162.610 52.600 162.910 ;
        RECT 62.220 162.870 62.820 163.170 ;
        RECT 63.420 162.870 64.920 163.170 ;
        RECT 65.520 162.870 66.120 163.170 ;
        RECT 31.245 162.335 34.445 162.425 ;
        RECT 30.655 161.915 34.445 162.335 ;
        RECT 46.600 162.010 48.100 162.610 ;
        RECT 51.400 162.010 52.900 162.610 ;
        RECT 62.220 162.570 62.520 162.870 ;
        RECT 61.920 162.270 62.520 162.570 ;
        RECT 30.655 161.795 33.840 161.915 ;
        RECT 30.070 161.395 33.840 161.795 ;
        RECT 46.900 161.710 48.700 162.010 ;
        RECT 50.800 161.710 52.600 162.010 ;
        RECT 61.920 161.970 62.820 162.270 ;
        RECT 63.720 161.970 64.620 162.870 ;
        RECT 65.820 162.570 66.120 162.870 ;
        RECT 77.370 163.130 78.270 163.430 ;
        RECT 79.170 163.130 80.070 164.030 ;
        RECT 81.270 163.730 81.570 164.030 ;
        RECT 93.980 163.880 95.480 164.480 ;
        RECT 81.270 163.430 81.870 163.730 ;
        RECT 93.380 163.580 94.580 163.880 ;
        RECT 94.880 163.580 96.080 163.880 ;
        RECT 80.970 163.130 81.870 163.430 ;
        RECT 91.880 163.280 93.980 163.580 ;
        RECT 95.480 163.280 97.880 163.580 ;
        RECT 65.820 162.270 66.420 162.570 ;
        RECT 65.520 161.970 66.420 162.270 ;
        RECT 47.800 161.410 49.000 161.710 ;
        RECT 50.500 161.410 51.700 161.710 ;
        RECT 30.070 161.245 33.245 161.395 ;
        RECT 29.495 160.870 33.245 161.245 ;
        RECT 48.400 161.110 49.600 161.410 ;
        RECT 49.900 161.110 51.100 161.410 ;
        RECT 29.495 160.690 32.655 160.870 ;
        RECT 28.925 160.335 32.655 160.690 ;
        RECT 49.000 160.510 50.500 161.110 ;
        RECT 61.920 160.770 66.420 161.970 ;
        RECT 77.370 161.930 81.870 163.130 ;
        RECT 91.580 162.980 93.380 163.280 ;
        RECT 96.080 162.980 97.880 163.280 ;
        RECT 91.580 162.680 92.780 162.980 ;
        RECT 96.680 162.680 97.880 162.980 ;
        RECT 91.580 162.380 92.480 162.680 ;
        RECT 96.980 162.380 97.880 162.680 ;
        RECT 91.880 162.080 92.180 162.380 ;
        RECT 93.680 162.080 93.980 162.380 ;
        RECT 94.280 162.080 94.580 162.380 ;
        RECT 94.880 162.080 95.180 162.380 ;
        RECT 95.480 162.080 95.780 162.380 ;
        RECT 97.280 162.080 97.580 162.380 ;
        RECT 104.630 162.260 105.080 168.740 ;
        RECT 105.345 168.675 109.385 168.740 ;
        RECT 105.345 168.345 110.055 168.675 ;
        RECT 106.030 168.235 110.055 168.345 ;
        RECT 106.030 167.940 110.720 168.235 ;
        RECT 106.715 167.785 110.720 167.940 ;
        RECT 106.715 167.525 111.380 167.785 ;
        RECT 107.385 167.330 111.380 167.525 ;
        RECT 107.385 167.105 112.035 167.330 ;
        RECT 108.055 166.865 112.035 167.105 ;
        RECT 108.055 166.675 112.680 166.865 ;
        RECT 108.720 166.395 112.680 166.675 ;
        RECT 108.720 166.235 113.320 166.395 ;
        RECT 109.380 165.915 113.320 166.235 ;
        RECT 109.380 165.785 113.955 165.915 ;
        RECT 110.035 165.425 113.955 165.785 ;
        RECT 110.035 165.330 114.585 165.425 ;
        RECT 110.680 164.930 114.585 165.330 ;
        RECT 110.680 164.865 115.210 164.930 ;
        RECT 111.320 164.425 115.210 164.865 ;
        RECT 111.320 164.395 115.825 164.425 ;
        RECT 111.955 163.915 115.825 164.395 ;
        RECT 112.585 163.425 116.435 163.915 ;
        RECT 113.210 163.395 116.435 163.425 ;
        RECT 107.110 163.030 109.510 163.330 ;
        RECT 106.810 162.730 109.510 163.030 ;
        RECT 113.210 162.930 117.040 163.395 ;
        RECT 113.825 162.870 117.040 162.930 ;
        RECT 106.210 162.130 110.110 162.730 ;
        RECT 113.825 162.425 117.635 162.870 ;
        RECT 114.435 162.335 117.635 162.425 ;
        RECT 28.925 160.125 32.070 160.335 ;
        RECT 48.400 160.210 49.600 160.510 ;
        RECT 49.900 160.210 51.100 160.510 ;
        RECT 28.360 159.795 32.070 160.125 ;
        RECT 46.900 159.910 49.000 160.210 ;
        RECT 50.500 159.910 52.900 160.210 ;
        RECT 28.360 159.555 31.495 159.795 ;
        RECT 27.805 159.245 31.495 159.555 ;
        RECT 46.600 159.610 48.400 159.910 ;
        RECT 51.100 159.610 52.900 159.910 ;
        RECT 46.600 159.310 47.800 159.610 ;
        RECT 51.700 159.310 52.900 159.610 ;
        RECT 27.805 158.980 30.925 159.245 ;
        RECT 46.600 159.010 47.500 159.310 ;
        RECT 52.000 159.010 52.900 159.310 ;
        RECT 60.640 159.180 61.200 160.570 ;
        RECT 62.220 160.170 66.120 160.770 ;
        RECT 76.090 160.340 76.650 161.730 ;
        RECT 77.670 161.330 81.570 161.930 ;
        RECT 93.680 161.480 95.780 162.080 ;
        RECT 78.270 161.030 80.970 161.330 ;
        RECT 93.380 161.180 94.280 161.480 ;
        RECT 95.180 161.180 96.380 161.480 ;
        RECT 78.570 160.730 80.970 161.030 ;
        RECT 92.780 160.880 94.580 161.180 ;
        RECT 94.880 160.880 96.380 161.180 ;
        RECT 105.910 160.930 110.410 162.130 ;
        RECT 114.435 161.915 118.225 162.335 ;
        RECT 115.040 161.795 118.225 161.915 ;
        RECT 115.040 161.395 118.810 161.795 ;
        RECT 92.780 160.580 93.380 160.880 ;
        RECT 93.980 160.580 95.480 160.880 ;
        RECT 96.080 160.580 96.680 160.880 ;
        RECT 62.820 159.870 65.520 160.170 ;
        RECT 63.120 159.570 65.520 159.870 ;
        RECT 27.255 158.970 30.925 158.980 ;
        RECT 27.255 158.520 34.550 158.970 ;
        RECT 46.900 158.710 47.200 159.010 ;
        RECT 48.700 158.710 49.000 159.010 ;
        RECT 49.300 158.710 49.600 159.010 ;
        RECT 49.900 158.710 50.200 159.010 ;
        RECT 50.500 158.710 50.800 159.010 ;
        RECT 52.300 158.710 52.600 159.010 ;
        RECT 27.255 158.395 30.360 158.520 ;
        RECT 26.715 158.125 30.360 158.395 ;
        RECT 26.715 157.805 29.805 158.125 ;
        RECT 26.180 157.555 29.805 157.805 ;
        RECT 26.180 157.210 29.255 157.555 ;
        RECT 25.655 156.980 29.255 157.210 ;
        RECT 25.655 156.605 28.715 156.980 ;
        RECT 34.100 156.970 34.550 158.520 ;
        RECT 48.700 158.110 50.800 158.710 ;
        RECT 36.580 157.740 38.980 158.040 ;
        RECT 48.400 157.810 49.300 158.110 ;
        RECT 50.200 157.810 51.400 158.110 ;
        RECT 36.280 157.440 38.980 157.740 ;
        RECT 47.800 157.510 49.600 157.810 ;
        RECT 49.900 157.510 51.400 157.810 ;
        RECT 35.680 156.840 39.580 157.440 ;
        RECT 47.800 157.210 48.400 157.510 ;
        RECT 49.000 157.210 50.500 157.510 ;
        RECT 51.100 157.210 51.700 157.510 ;
        RECT 47.800 156.910 48.100 157.210 ;
        RECT 25.135 156.395 28.715 156.605 ;
        RECT 25.135 155.995 28.180 156.395 ;
        RECT 24.625 155.805 28.180 155.995 ;
        RECT 24.625 155.380 27.655 155.805 ;
        RECT 24.120 155.210 27.655 155.380 ;
        RECT 35.380 155.640 39.880 156.840 ;
        RECT 35.380 155.340 36.280 155.640 ;
        RECT 24.120 154.755 27.135 155.210 ;
        RECT 35.380 155.040 35.980 155.340 ;
        RECT 23.625 154.605 27.135 154.755 ;
        RECT 35.680 154.740 35.980 155.040 ;
        RECT 37.180 154.740 38.080 155.640 ;
        RECT 38.980 155.340 39.880 155.640 ;
        RECT 39.280 155.040 39.880 155.340 ;
        RECT 47.500 156.610 48.100 156.910 ;
        RECT 47.500 156.310 48.400 156.610 ;
        RECT 49.300 156.310 50.200 157.210 ;
        RECT 51.400 156.910 51.700 157.210 ;
        RECT 51.400 156.610 52.000 156.910 ;
        RECT 51.100 156.310 52.000 156.610 ;
        RECT 47.500 155.110 52.000 156.310 ;
        RECT 60.640 155.905 61.090 159.180 ;
        RECT 73.445 157.600 75.440 157.610 ;
        RECT 76.090 157.600 76.540 160.340 ;
        RECT 92.780 160.280 93.080 160.580 ;
        RECT 92.480 159.980 93.080 160.280 ;
        RECT 92.480 159.680 93.380 159.980 ;
        RECT 94.280 159.680 95.180 160.580 ;
        RECT 96.380 160.280 96.680 160.580 ;
        RECT 105.910 160.630 106.810 160.930 ;
        RECT 105.910 160.330 106.510 160.630 ;
        RECT 96.380 159.980 96.980 160.280 ;
        RECT 96.080 159.680 96.980 159.980 ;
        RECT 92.480 158.480 96.980 159.680 ;
        RECT 106.210 160.030 106.510 160.330 ;
        RECT 107.710 160.030 108.610 160.930 ;
        RECT 109.510 160.630 110.410 160.930 ;
        RECT 115.635 161.245 118.810 161.395 ;
        RECT 115.635 160.870 119.385 161.245 ;
        RECT 109.810 160.330 110.410 160.630 ;
        RECT 116.225 160.690 119.385 160.870 ;
        RECT 116.225 160.335 119.955 160.690 ;
        RECT 109.810 160.030 110.110 160.330 ;
        RECT 106.210 159.730 106.810 160.030 ;
        RECT 107.410 159.730 108.910 160.030 ;
        RECT 109.510 159.730 110.110 160.030 ;
        RECT 116.810 160.125 119.955 160.335 ;
        RECT 116.810 159.795 120.520 160.125 ;
        RECT 106.210 159.430 108.010 159.730 ;
        RECT 108.310 159.430 109.810 159.730 ;
        RECT 106.810 159.130 107.710 159.430 ;
        RECT 108.610 159.130 109.810 159.430 ;
        RECT 117.385 159.555 120.520 159.795 ;
        RECT 117.385 159.245 121.075 159.555 ;
        RECT 107.110 158.530 109.210 159.130 ;
        RECT 117.955 158.980 121.075 159.245 ;
        RECT 117.955 158.690 121.625 158.980 ;
        RECT 72.710 157.580 76.540 157.600 ;
        RECT 71.975 157.550 76.905 157.580 ;
        RECT 71.245 157.505 77.635 157.550 ;
        RECT 70.515 157.450 78.365 157.505 ;
        RECT 69.780 157.375 79.100 157.450 ;
        RECT 69.050 157.295 79.830 157.375 ;
        RECT 68.325 157.200 80.555 157.295 ;
        RECT 67.595 157.090 81.285 157.200 ;
        RECT 66.870 156.970 82.010 157.090 ;
        RECT 66.150 156.835 82.730 156.970 ;
        RECT 91.200 156.890 91.760 158.280 ;
        RECT 92.780 157.880 96.680 158.480 ;
        RECT 105.310 158.230 106.210 158.530 ;
        RECT 107.110 158.230 107.410 158.530 ;
        RECT 107.710 158.230 108.010 158.530 ;
        RECT 108.310 158.230 108.610 158.530 ;
        RECT 108.910 158.230 109.210 158.530 ;
        RECT 110.110 158.230 111.010 158.530 ;
        RECT 118.520 158.395 121.625 158.690 ;
        RECT 93.380 157.580 96.080 157.880 ;
        RECT 105.010 157.630 106.510 158.230 ;
        RECT 109.810 157.630 111.310 158.230 ;
        RECT 118.520 158.125 122.165 158.395 ;
        RECT 119.075 157.805 122.165 158.125 ;
        RECT 93.680 157.280 96.080 157.580 ;
        RECT 105.310 157.330 107.110 157.630 ;
        RECT 109.210 157.330 111.010 157.630 ;
        RECT 119.075 157.555 122.700 157.805 ;
        RECT 106.210 157.030 107.410 157.330 ;
        RECT 108.910 157.030 110.110 157.330 ;
        RECT 119.625 157.210 122.700 157.555 ;
        RECT 65.430 156.690 83.450 156.835 ;
        RECT 64.710 156.530 84.170 156.690 ;
        RECT 63.995 156.360 84.885 156.530 ;
        RECT 63.280 156.175 85.600 156.360 ;
        RECT 62.570 155.980 86.310 156.175 ;
        RECT 60.640 155.770 61.345 155.905 ;
        RECT 61.865 155.770 87.015 155.980 ;
        RECT 60.640 155.600 87.715 155.770 ;
        RECT 60.640 155.580 73.975 155.600 ;
        RECT 74.905 155.580 87.715 155.600 ;
        RECT 60.640 155.550 73.245 155.580 ;
        RECT 75.635 155.550 87.715 155.580 ;
        RECT 60.465 155.505 72.515 155.550 ;
        RECT 76.365 155.505 88.415 155.550 ;
        RECT 60.465 155.450 71.780 155.505 ;
        RECT 77.100 155.450 88.415 155.505 ;
        RECT 60.465 155.375 71.050 155.450 ;
        RECT 77.830 155.375 88.415 155.450 ;
        RECT 60.465 155.320 70.325 155.375 ;
        RECT 59.770 155.295 70.325 155.320 ;
        RECT 78.555 155.320 88.415 155.375 ;
        RECT 78.555 155.295 89.110 155.320 ;
        RECT 59.770 155.200 69.595 155.295 ;
        RECT 79.285 155.200 89.110 155.295 ;
        RECT 39.280 154.740 39.580 155.040 ;
        RECT 23.625 154.125 26.625 154.605 ;
        RECT 35.680 154.440 36.280 154.740 ;
        RECT 36.880 154.440 38.380 154.740 ;
        RECT 38.980 154.440 39.580 154.740 ;
        RECT 35.680 154.140 37.480 154.440 ;
        RECT 37.780 154.140 39.280 154.440 ;
        RECT 23.135 153.995 26.625 154.125 ;
        RECT 23.135 153.490 26.120 153.995 ;
        RECT 36.280 153.840 37.180 154.140 ;
        RECT 38.080 153.840 39.280 154.140 ;
        RECT 22.655 153.380 26.120 153.490 ;
        RECT 22.655 152.850 25.625 153.380 ;
        RECT 36.580 153.240 38.680 153.840 ;
        RECT 46.220 153.520 46.780 154.910 ;
        RECT 47.800 154.510 51.700 155.110 ;
        RECT 59.770 155.090 68.870 155.200 ;
        RECT 80.010 155.090 89.110 155.200 ;
        RECT 59.770 155.075 68.150 155.090 ;
        RECT 59.080 154.970 68.150 155.075 ;
        RECT 80.730 155.075 89.110 155.090 ;
        RECT 80.730 154.970 89.800 155.075 ;
        RECT 59.080 154.835 67.430 154.970 ;
        RECT 81.450 154.835 89.800 154.970 ;
        RECT 59.080 154.820 66.710 154.835 ;
        RECT 58.390 154.690 66.710 154.820 ;
        RECT 82.170 154.820 89.800 154.835 ;
        RECT 82.170 154.690 90.490 154.820 ;
        RECT 58.390 154.550 65.995 154.690 ;
        RECT 57.710 154.530 65.995 154.550 ;
        RECT 82.885 154.550 90.490 154.690 ;
        RECT 91.200 154.635 91.650 156.890 ;
        RECT 106.810 156.730 108.010 157.030 ;
        RECT 108.310 156.730 109.510 157.030 ;
        RECT 119.625 156.980 123.225 157.210 ;
        RECT 107.410 156.130 108.910 156.730 ;
        RECT 120.165 156.605 123.225 156.980 ;
        RECT 120.165 156.395 123.745 156.605 ;
        RECT 106.810 155.830 108.010 156.130 ;
        RECT 108.310 155.830 109.510 156.130 ;
        RECT 120.700 155.995 123.745 156.395 ;
        RECT 105.310 155.530 107.410 155.830 ;
        RECT 108.910 155.530 111.310 155.830 ;
        RECT 120.700 155.805 124.255 155.995 ;
        RECT 90.865 154.550 91.650 154.635 ;
        RECT 105.010 155.230 106.810 155.530 ;
        RECT 109.510 155.230 111.310 155.530 ;
        RECT 105.010 154.930 106.210 155.230 ;
        RECT 110.110 154.930 111.310 155.230 ;
        RECT 121.225 155.380 124.255 155.805 ;
        RECT 121.225 155.210 124.760 155.380 ;
        RECT 105.010 154.630 105.910 154.930 ;
        RECT 110.410 154.630 111.310 154.930 ;
        RECT 121.745 154.755 124.760 155.210 ;
        RECT 121.745 154.635 125.255 154.755 ;
        RECT 82.885 154.530 91.650 154.550 ;
        RECT 48.400 154.210 51.100 154.510 ;
        RECT 57.710 154.360 65.280 154.530 ;
        RECT 83.600 154.360 91.650 154.530 ;
        RECT 57.710 154.270 64.570 154.360 ;
        RECT 48.700 153.910 51.100 154.210 ;
        RECT 57.030 154.175 64.570 154.270 ;
        RECT 84.310 154.270 91.650 154.360 ;
        RECT 105.310 154.330 105.610 154.630 ;
        RECT 107.110 154.330 107.410 154.630 ;
        RECT 107.710 154.330 108.010 154.630 ;
        RECT 108.310 154.330 108.610 154.630 ;
        RECT 108.910 154.330 109.210 154.630 ;
        RECT 110.710 154.330 111.010 154.630 ;
        RECT 84.310 154.175 91.850 154.270 ;
        RECT 57.030 153.980 63.865 154.175 ;
        RECT 85.015 153.980 91.850 154.175 ;
        RECT 57.030 153.975 63.165 153.980 ;
        RECT 56.360 153.770 63.165 153.975 ;
        RECT 85.715 153.975 91.850 153.980 ;
        RECT 85.715 153.770 92.520 153.975 ;
        RECT 56.360 153.670 62.465 153.770 ;
        RECT 55.695 153.550 62.465 153.670 ;
        RECT 86.415 153.670 92.520 153.770 ;
        RECT 107.110 153.730 109.210 154.330 ;
        RECT 115.170 154.185 125.255 154.635 ;
        RECT 86.415 153.550 93.185 153.670 ;
        RECT 34.780 152.940 35.680 153.240 ;
        RECT 36.580 152.940 36.880 153.240 ;
        RECT 37.180 152.940 37.480 153.240 ;
        RECT 37.780 152.940 38.080 153.240 ;
        RECT 38.380 152.940 38.680 153.240 ;
        RECT 39.580 152.940 40.480 153.240 ;
        RECT 22.185 152.755 25.625 152.850 ;
        RECT 22.185 152.205 25.135 152.755 ;
        RECT 34.480 152.340 35.980 152.940 ;
        RECT 39.280 152.340 40.780 152.940 ;
        RECT 21.720 152.125 25.135 152.205 ;
        RECT 21.720 151.550 24.655 152.125 ;
        RECT 34.780 152.040 36.580 152.340 ;
        RECT 38.680 152.040 40.480 152.340 ;
        RECT 35.680 151.740 36.880 152.040 ;
        RECT 38.380 151.740 39.580 152.040 ;
        RECT 21.265 151.490 24.655 151.550 ;
        RECT 21.265 150.890 24.185 151.490 ;
        RECT 36.280 151.440 37.480 151.740 ;
        RECT 37.780 151.440 38.980 151.740 ;
        RECT 20.815 150.850 24.185 150.890 ;
        RECT 20.815 150.225 23.720 150.850 ;
        RECT 36.880 150.840 38.380 151.440 ;
        RECT 36.280 150.540 37.480 150.840 ;
        RECT 37.780 150.540 38.980 150.840 ;
        RECT 34.780 150.240 36.880 150.540 ;
        RECT 38.380 150.240 40.780 150.540 ;
        RECT 20.375 150.205 23.720 150.225 ;
        RECT 20.375 149.555 23.265 150.205 ;
        RECT 19.945 149.550 23.265 149.555 ;
        RECT 34.480 149.940 36.280 150.240 ;
        RECT 38.980 149.940 40.780 150.240 ;
        RECT 34.480 149.640 35.680 149.940 ;
        RECT 39.580 149.640 40.780 149.940 ;
        RECT 19.945 148.890 22.815 149.550 ;
        RECT 34.480 149.340 35.380 149.640 ;
        RECT 39.880 149.340 40.780 149.640 ;
        RECT 34.780 149.040 35.080 149.340 ;
        RECT 36.580 149.040 36.880 149.340 ;
        RECT 37.180 149.040 37.480 149.340 ;
        RECT 37.780 149.040 38.080 149.340 ;
        RECT 38.380 149.040 38.680 149.340 ;
        RECT 40.180 149.040 40.480 149.340 ;
        RECT 19.945 148.885 22.375 148.890 ;
        RECT 19.525 148.225 22.375 148.885 ;
        RECT 36.580 148.440 38.680 149.040 ;
        RECT 19.525 148.200 21.945 148.225 ;
        RECT 19.110 147.835 21.945 148.200 ;
        RECT 36.280 148.140 37.180 148.440 ;
        RECT 38.080 148.140 39.280 148.440 ;
        RECT 35.680 147.840 37.480 148.140 ;
        RECT 37.780 147.840 39.280 148.140 ;
        RECT 19.110 147.515 25.810 147.835 ;
        RECT 18.705 147.385 25.810 147.515 ;
        RECT 18.705 146.885 21.525 147.385 ;
        RECT 18.705 146.825 21.110 146.885 ;
        RECT 18.310 146.200 21.110 146.825 ;
        RECT 18.310 146.130 20.705 146.200 ;
        RECT 25.360 146.170 25.810 147.385 ;
        RECT 35.680 147.540 36.280 147.840 ;
        RECT 36.880 147.540 38.380 147.840 ;
        RECT 38.980 147.540 39.580 147.840 ;
        RECT 35.680 147.240 35.980 147.540 ;
        RECT 27.840 146.940 30.240 147.240 ;
        RECT 27.540 146.640 30.240 146.940 ;
        RECT 35.380 146.940 35.980 147.240 ;
        RECT 35.380 146.640 36.280 146.940 ;
        RECT 37.180 146.640 38.080 147.540 ;
        RECT 39.280 147.240 39.580 147.540 ;
        RECT 46.220 147.780 46.670 153.520 ;
        RECT 55.695 153.355 61.770 153.550 ;
        RECT 55.030 153.320 61.770 153.355 ;
        RECT 87.110 153.355 93.185 153.550 ;
        RECT 106.810 153.430 107.710 153.730 ;
        RECT 108.610 153.430 109.810 153.730 ;
        RECT 87.110 153.320 93.850 153.355 ;
        RECT 55.030 153.075 61.080 153.320 ;
        RECT 87.800 153.075 93.850 153.320 ;
        RECT 55.030 153.030 60.390 153.075 ;
        RECT 54.375 152.820 60.390 153.030 ;
        RECT 88.490 153.030 93.850 153.075 ;
        RECT 106.210 153.130 108.010 153.430 ;
        RECT 108.310 153.130 109.810 153.430 ;
        RECT 88.490 152.820 94.505 153.030 ;
        RECT 54.375 152.690 59.710 152.820 ;
        RECT 53.725 152.550 59.710 152.690 ;
        RECT 89.170 152.690 94.505 152.820 ;
        RECT 106.210 152.830 106.810 153.130 ;
        RECT 107.410 152.830 108.910 153.130 ;
        RECT 109.510 152.830 110.110 153.130 ;
        RECT 89.170 152.550 95.155 152.690 ;
        RECT 53.725 152.340 59.030 152.550 ;
        RECT 53.080 152.270 59.030 152.340 ;
        RECT 89.850 152.340 95.155 152.550 ;
        RECT 106.210 152.530 106.510 152.830 ;
        RECT 89.850 152.270 95.800 152.340 ;
        RECT 53.080 151.980 58.360 152.270 ;
        RECT 52.445 151.975 58.360 151.980 ;
        RECT 90.520 151.980 95.800 152.270 ;
        RECT 105.910 152.230 106.510 152.530 ;
        RECT 90.520 151.975 96.440 151.980 ;
        RECT 52.445 151.670 57.695 151.975 ;
        RECT 91.185 151.670 96.440 151.975 ;
        RECT 52.445 151.610 57.030 151.670 ;
        RECT 51.810 151.355 57.030 151.610 ;
        RECT 91.850 151.610 96.440 151.670 ;
        RECT 105.910 151.930 106.810 152.230 ;
        RECT 107.710 151.930 108.610 152.830 ;
        RECT 109.810 152.530 110.110 152.830 ;
        RECT 109.810 152.230 110.410 152.530 ;
        RECT 109.510 151.930 110.410 152.230 ;
        RECT 91.850 151.355 97.070 151.610 ;
        RECT 51.810 151.225 56.375 151.355 ;
        RECT 51.185 151.030 56.375 151.225 ;
        RECT 92.505 151.225 97.070 151.355 ;
        RECT 92.505 151.030 97.695 151.225 ;
        RECT 51.185 150.830 55.725 151.030 ;
        RECT 50.570 150.690 55.725 150.830 ;
        RECT 93.155 150.830 97.695 151.030 ;
        RECT 93.155 150.690 98.310 150.830 ;
        RECT 105.910 150.730 110.410 151.930 ;
        RECT 115.170 150.900 115.620 154.185 ;
        RECT 122.255 154.125 125.255 154.185 ;
        RECT 122.255 153.995 125.745 154.125 ;
        RECT 122.760 153.490 125.745 153.995 ;
        RECT 122.760 153.380 126.225 153.490 ;
        RECT 123.255 152.850 126.225 153.380 ;
        RECT 123.255 152.755 126.695 152.850 ;
        RECT 123.745 152.205 126.695 152.755 ;
        RECT 123.745 152.125 127.160 152.205 ;
        RECT 117.650 151.670 120.050 151.970 ;
        RECT 117.350 151.370 120.050 151.670 ;
        RECT 124.225 151.550 127.160 152.125 ;
        RECT 124.225 151.490 127.615 151.550 ;
        RECT 116.750 150.770 120.650 151.370 ;
        RECT 124.695 150.890 127.615 151.490 ;
        RECT 124.695 150.850 128.065 150.890 ;
        RECT 50.570 150.425 55.080 150.690 ;
        RECT 49.955 150.340 55.080 150.425 ;
        RECT 49.955 150.010 54.445 150.340 ;
        RECT 49.350 149.980 54.445 150.010 ;
        RECT 49.350 149.610 53.810 149.980 ;
        RECT 49.350 149.585 53.185 149.610 ;
        RECT 48.755 149.225 53.185 149.585 ;
        RECT 48.755 149.150 52.570 149.225 ;
        RECT 48.165 148.830 52.570 149.150 ;
        RECT 48.165 148.705 51.955 148.830 ;
        RECT 47.585 148.425 51.955 148.705 ;
        RECT 47.585 148.250 51.350 148.425 ;
        RECT 66.380 148.410 84.060 150.620 ;
        RECT 93.800 150.425 98.310 150.690 ;
        RECT 93.800 150.340 98.925 150.425 ;
        RECT 94.440 150.010 98.925 150.340 ;
        RECT 94.440 149.980 99.530 150.010 ;
        RECT 95.070 149.610 99.530 149.980 ;
        RECT 95.695 149.585 99.530 149.610 ;
        RECT 95.695 149.225 100.125 149.585 ;
        RECT 96.310 149.150 100.125 149.225 ;
        RECT 96.310 148.830 100.715 149.150 ;
        RECT 96.925 148.705 100.715 148.830 ;
        RECT 104.630 149.140 105.190 150.530 ;
        RECT 106.210 150.130 110.110 150.730 ;
        RECT 106.810 149.830 109.510 150.130 ;
        RECT 107.110 149.530 109.510 149.830 ;
        RECT 116.450 149.570 120.950 150.770 ;
        RECT 125.160 150.225 128.065 150.850 ;
        RECT 125.160 150.205 128.505 150.225 ;
        RECT 116.450 149.270 117.350 149.570 ;
        RECT 96.925 148.475 101.295 148.705 ;
        RECT 104.630 148.475 105.080 149.140 ;
        RECT 116.450 148.970 117.050 149.270 ;
        RECT 96.925 148.425 105.080 148.475 ;
        RECT 47.010 148.010 51.350 148.250 ;
        RECT 47.010 147.780 50.755 148.010 ;
        RECT 46.220 147.585 50.755 147.780 ;
        RECT 46.220 147.305 50.165 147.585 ;
        RECT 39.280 146.940 39.880 147.240 ;
        RECT 38.980 146.640 39.880 146.940 ;
        RECT 45.890 147.150 50.165 147.305 ;
        RECT 45.890 146.820 49.585 147.150 ;
        RECT 17.920 145.515 20.705 146.130 ;
        RECT 26.940 146.040 30.840 146.640 ;
        RECT 17.920 145.430 20.310 145.515 ;
        RECT 17.540 144.825 20.310 145.430 ;
        RECT 26.640 144.840 31.140 146.040 ;
        RECT 35.380 145.440 39.880 146.640 ;
        RECT 45.340 146.705 49.585 146.820 ;
        RECT 45.340 146.325 49.010 146.705 ;
        RECT 44.800 146.250 49.010 146.325 ;
        RECT 44.800 145.820 48.445 146.250 ;
        RECT 64.170 146.200 84.060 148.410 ;
        RECT 97.530 148.025 105.080 148.425 ;
        RECT 116.750 148.670 117.050 148.970 ;
        RECT 118.250 148.670 119.150 149.570 ;
        RECT 120.050 149.270 120.950 149.570 ;
        RECT 125.615 149.555 128.505 150.205 ;
        RECT 125.615 149.550 128.935 149.555 ;
        RECT 120.350 148.970 120.950 149.270 ;
        RECT 120.350 148.670 120.650 148.970 ;
        RECT 126.065 148.890 128.935 149.550 ;
        RECT 116.750 148.370 117.350 148.670 ;
        RECT 117.950 148.370 119.450 148.670 ;
        RECT 120.050 148.370 120.650 148.670 ;
        RECT 126.505 148.885 128.935 148.890 ;
        RECT 116.750 148.070 118.550 148.370 ;
        RECT 118.850 148.070 120.350 148.370 ;
        RECT 126.505 148.225 129.355 148.885 ;
        RECT 97.530 148.010 101.870 148.025 ;
        RECT 98.125 147.780 101.870 148.010 ;
        RECT 98.125 147.585 102.435 147.780 ;
        RECT 117.350 147.770 118.250 148.070 ;
        RECT 119.150 147.770 120.350 148.070 ;
        RECT 126.935 148.200 129.355 148.225 ;
        RECT 98.715 147.305 102.435 147.585 ;
        RECT 98.715 147.150 102.990 147.305 ;
        RECT 117.650 147.170 119.750 147.770 ;
        RECT 126.935 147.555 129.770 148.200 ;
        RECT 127.355 147.515 129.770 147.555 ;
        RECT 99.295 146.820 102.990 147.150 ;
        RECT 115.850 146.870 116.750 147.170 ;
        RECT 117.650 146.870 117.950 147.170 ;
        RECT 118.250 146.870 118.550 147.170 ;
        RECT 118.850 146.870 119.150 147.170 ;
        RECT 119.450 146.870 119.750 147.170 ;
        RECT 120.650 146.870 121.550 147.170 ;
        RECT 127.355 146.885 130.175 147.515 ;
        RECT 99.295 146.705 103.540 146.820 ;
        RECT 99.870 146.325 103.540 146.705 ;
        RECT 99.870 146.250 104.080 146.325 ;
        RECT 115.550 146.270 117.050 146.870 ;
        RECT 120.350 146.270 121.850 146.870 ;
        RECT 127.770 146.825 130.175 146.885 ;
        RECT 44.265 145.780 48.445 145.820 ;
        RECT 17.540 144.725 19.920 144.825 ;
        RECT 17.170 144.130 19.920 144.725 ;
        RECT 26.640 144.540 27.540 144.840 ;
        RECT 26.640 144.240 27.240 144.540 ;
        RECT 17.170 144.015 19.540 144.130 ;
        RECT 16.810 143.430 19.540 144.015 ;
        RECT 26.940 143.940 27.240 144.240 ;
        RECT 28.440 143.940 29.340 144.840 ;
        RECT 30.240 144.540 31.140 144.840 ;
        RECT 30.540 144.240 31.140 144.540 ;
        RECT 30.540 143.940 30.840 144.240 ;
        RECT 26.940 143.640 27.540 143.940 ;
        RECT 28.140 143.640 29.640 143.940 ;
        RECT 30.240 143.640 30.840 143.940 ;
        RECT 34.100 143.850 34.660 145.240 ;
        RECT 35.680 144.840 39.580 145.440 ;
        RECT 44.265 145.305 47.890 145.780 ;
        RECT 36.280 144.540 38.980 144.840 ;
        RECT 43.745 144.820 47.340 145.305 ;
        RECT 43.745 144.785 46.800 144.820 ;
        RECT 36.580 144.240 38.980 144.540 ;
        RECT 43.230 144.325 46.800 144.785 ;
        RECT 43.230 144.250 46.265 144.325 ;
        RECT 16.810 143.305 19.170 143.430 ;
        RECT 26.940 143.340 28.740 143.640 ;
        RECT 29.040 143.340 30.540 143.640 ;
        RECT 16.455 142.725 19.170 143.305 ;
        RECT 27.540 143.040 28.440 143.340 ;
        RECT 29.340 143.040 30.540 143.340 ;
        RECT 34.100 143.435 34.550 143.850 ;
        RECT 42.725 143.820 46.265 144.250 ;
        RECT 42.725 143.710 45.745 143.820 ;
        RECT 42.230 143.435 45.745 143.710 ;
        RECT 34.100 143.305 45.745 143.435 ;
        RECT 16.455 142.585 18.810 142.725 ;
        RECT 16.115 142.015 18.810 142.585 ;
        RECT 27.840 142.440 29.940 143.040 ;
        RECT 34.100 142.985 45.230 143.305 ;
        RECT 34.100 142.970 34.550 142.985 ;
        RECT 41.745 142.785 45.230 142.985 ;
        RECT 41.745 142.605 44.725 142.785 ;
        RECT 26.040 142.140 26.940 142.440 ;
        RECT 27.840 142.140 28.140 142.440 ;
        RECT 28.440 142.140 28.740 142.440 ;
        RECT 29.040 142.140 29.340 142.440 ;
        RECT 29.640 142.140 29.940 142.440 ;
        RECT 30.840 142.140 31.740 142.440 ;
        RECT 41.270 142.250 44.725 142.605 ;
        RECT 16.115 141.860 18.455 142.015 ;
        RECT 15.780 141.305 18.455 141.860 ;
        RECT 25.740 141.540 27.240 142.140 ;
        RECT 30.540 141.540 32.040 142.140 ;
        RECT 41.270 142.040 44.230 142.250 ;
        RECT 40.800 141.710 44.230 142.040 ;
        RECT 59.750 141.780 88.480 146.200 ;
        RECT 100.435 145.820 104.080 146.250 ;
        RECT 115.850 145.970 117.650 146.270 ;
        RECT 119.750 145.970 121.550 146.270 ;
        RECT 127.770 146.200 130.570 146.825 ;
        RECT 128.175 146.130 130.570 146.200 ;
        RECT 100.435 145.780 104.615 145.820 ;
        RECT 100.990 145.305 104.615 145.780 ;
        RECT 116.750 145.670 117.950 145.970 ;
        RECT 119.450 145.670 120.650 145.970 ;
        RECT 117.350 145.370 118.550 145.670 ;
        RECT 118.850 145.370 120.050 145.670 ;
        RECT 128.175 145.515 130.960 146.130 ;
        RECT 128.570 145.430 130.960 145.515 ;
        RECT 101.540 144.820 105.135 145.305 ;
        RECT 102.080 144.785 105.135 144.820 ;
        RECT 102.080 144.325 105.650 144.785 ;
        RECT 117.950 144.770 119.450 145.370 ;
        RECT 128.570 144.825 131.340 145.430 ;
        RECT 117.350 144.470 118.550 144.770 ;
        RECT 118.850 144.470 120.050 144.770 ;
        RECT 128.960 144.725 131.340 144.825 ;
        RECT 102.615 144.250 105.650 144.325 ;
        RECT 102.615 143.820 106.155 144.250 ;
        RECT 115.850 144.170 117.950 144.470 ;
        RECT 119.450 144.170 121.850 144.470 ;
        RECT 103.135 143.710 106.155 143.820 ;
        RECT 115.550 143.870 117.350 144.170 ;
        RECT 120.050 143.870 121.850 144.170 ;
        RECT 128.960 144.130 131.710 144.725 ;
        RECT 103.135 143.305 106.650 143.710 ;
        RECT 103.650 143.160 106.650 143.305 ;
        RECT 115.550 143.570 116.750 143.870 ;
        RECT 120.650 143.570 121.850 143.870 ;
        RECT 115.550 143.270 116.450 143.570 ;
        RECT 120.950 143.270 121.850 143.570 ;
        RECT 129.340 144.015 131.710 144.130 ;
        RECT 129.340 143.430 132.070 144.015 ;
        RECT 129.710 143.305 132.070 143.430 ;
        RECT 103.650 142.785 107.135 143.160 ;
        RECT 115.850 142.970 116.150 143.270 ;
        RECT 117.650 142.970 117.950 143.270 ;
        RECT 118.250 142.970 118.550 143.270 ;
        RECT 118.850 142.970 119.150 143.270 ;
        RECT 119.450 142.970 119.750 143.270 ;
        RECT 121.250 142.970 121.550 143.270 ;
        RECT 104.155 142.605 107.135 142.785 ;
        RECT 104.155 142.250 107.610 142.605 ;
        RECT 117.650 142.370 119.750 142.970 ;
        RECT 129.710 142.725 132.425 143.305 ;
        RECT 130.070 142.585 132.425 142.725 ;
        RECT 104.650 142.040 107.610 142.250 ;
        RECT 117.350 142.070 118.250 142.370 ;
        RECT 119.150 142.070 120.350 142.370 ;
        RECT 15.780 141.135 18.115 141.305 ;
        RECT 26.040 141.240 27.840 141.540 ;
        RECT 29.940 141.240 31.740 141.540 ;
        RECT 40.800 141.465 43.745 141.710 ;
        RECT 15.455 140.585 18.115 141.135 ;
        RECT 26.940 140.940 28.140 141.240 ;
        RECT 29.640 140.940 30.840 141.240 ;
        RECT 40.345 141.160 43.745 141.465 ;
        RECT 27.540 140.640 28.740 140.940 ;
        RECT 29.040 140.640 30.240 140.940 ;
        RECT 40.345 140.885 43.270 141.160 ;
        RECT 15.455 140.405 17.780 140.585 ;
        RECT 15.135 139.860 17.780 140.405 ;
        RECT 28.140 140.040 29.640 140.640 ;
        RECT 39.900 140.605 43.270 140.885 ;
        RECT 39.900 140.295 42.800 140.605 ;
        RECT 39.465 140.040 42.800 140.295 ;
        RECT 15.135 139.670 17.455 139.860 ;
        RECT 27.540 139.740 28.740 140.040 ;
        RECT 29.040 139.740 30.240 140.040 ;
        RECT 14.830 139.135 17.455 139.670 ;
        RECT 26.040 139.440 28.140 139.740 ;
        RECT 29.640 139.440 32.040 139.740 ;
        RECT 39.465 139.700 42.345 140.040 ;
        RECT 25.740 139.140 27.540 139.440 ;
        RECT 30.240 139.140 32.040 139.440 ;
        RECT 14.830 138.930 17.135 139.135 ;
        RECT 14.530 138.405 17.135 138.930 ;
        RECT 25.740 138.840 26.940 139.140 ;
        RECT 30.840 138.840 32.040 139.140 ;
        RECT 39.040 139.465 42.345 139.700 ;
        RECT 39.040 139.095 41.900 139.465 ;
        RECT 25.740 138.540 26.640 138.840 ;
        RECT 31.140 138.540 32.040 138.840 ;
        RECT 38.625 138.885 41.900 139.095 ;
        RECT 14.530 138.190 16.830 138.405 ;
        RECT 26.040 138.240 26.340 138.540 ;
        RECT 27.840 138.240 28.140 138.540 ;
        RECT 28.440 138.240 28.740 138.540 ;
        RECT 29.040 138.240 29.340 138.540 ;
        RECT 29.640 138.240 29.940 138.540 ;
        RECT 31.440 138.240 31.740 138.540 ;
        RECT 38.625 138.480 41.465 138.885 ;
        RECT 38.220 138.295 41.465 138.480 ;
        RECT 14.245 137.670 16.830 138.190 ;
        RECT 14.245 137.445 16.530 137.670 ;
        RECT 27.840 137.640 29.940 138.240 ;
        RECT 38.220 137.865 41.040 138.295 ;
        RECT 37.825 137.700 41.040 137.865 ;
        RECT 13.965 136.930 16.530 137.445 ;
        RECT 27.540 137.340 28.440 137.640 ;
        RECT 29.340 137.340 30.540 137.640 ;
        RECT 26.940 137.040 28.740 137.340 ;
        RECT 29.040 137.040 30.540 137.340 ;
        RECT 37.825 137.240 40.625 137.700 ;
        RECT 37.440 137.095 40.625 137.240 ;
        RECT 13.965 136.695 16.245 136.930 ;
        RECT 13.695 136.190 16.245 136.695 ;
        RECT 26.940 136.740 27.540 137.040 ;
        RECT 28.140 136.740 29.640 137.040 ;
        RECT 30.240 136.740 30.840 137.040 ;
        RECT 26.940 136.440 27.240 136.740 ;
        RECT 13.695 135.940 15.965 136.190 ;
        RECT 13.435 135.445 15.965 135.940 ;
        RECT 26.640 136.140 27.240 136.440 ;
        RECT 26.640 135.840 27.540 136.140 ;
        RECT 28.440 135.840 29.340 136.740 ;
        RECT 30.540 136.440 30.840 136.740 ;
        RECT 37.440 136.605 40.220 137.095 ;
        RECT 37.070 136.480 40.220 136.605 ;
        RECT 30.540 136.140 31.140 136.440 ;
        RECT 30.240 135.840 31.140 136.140 ;
        RECT 37.070 135.970 39.825 136.480 ;
        RECT 13.435 135.185 15.695 135.445 ;
        RECT 13.185 134.695 15.695 135.185 ;
        RECT 13.185 134.430 15.435 134.695 ;
        RECT 26.640 134.640 31.140 135.840 ;
        RECT 36.710 135.865 39.825 135.970 ;
        RECT 36.710 135.325 39.440 135.865 ;
        RECT 36.360 135.240 39.440 135.325 ;
        RECT 36.360 134.675 39.070 135.240 ;
        RECT 12.940 133.940 15.435 134.430 ;
        RECT 12.940 133.665 15.185 133.940 ;
        RECT 12.710 133.185 15.185 133.665 ;
        RECT 12.710 132.900 14.940 133.185 ;
        RECT 12.490 132.430 14.940 132.900 ;
        RECT 25.360 133.050 25.920 134.440 ;
        RECT 26.940 134.040 30.840 134.640 ;
        RECT 36.020 134.605 39.070 134.675 ;
        RECT 27.540 133.740 30.240 134.040 ;
        RECT 36.020 134.020 38.710 134.605 ;
        RECT 27.840 133.440 30.240 133.740 ;
        RECT 35.695 133.970 38.710 134.020 ;
        RECT 35.695 133.355 38.360 133.970 ;
        RECT 35.380 133.325 38.360 133.355 ;
        RECT 25.360 132.620 25.810 133.050 ;
        RECT 35.380 132.690 38.020 133.325 ;
        RECT 35.075 132.675 38.020 132.690 ;
        RECT 57.540 132.940 90.690 141.780 ;
        RECT 104.650 141.710 108.080 142.040 ;
        RECT 105.135 141.465 108.080 141.710 ;
        RECT 116.750 141.770 118.550 142.070 ;
        RECT 118.850 141.770 120.350 142.070 ;
        RECT 130.070 142.015 132.765 142.585 ;
        RECT 130.425 141.860 132.765 142.015 ;
        RECT 116.750 141.470 117.350 141.770 ;
        RECT 117.950 141.470 119.450 141.770 ;
        RECT 120.050 141.470 120.650 141.770 ;
        RECT 105.135 141.160 108.535 141.465 ;
        RECT 116.750 141.170 117.050 141.470 ;
        RECT 105.610 140.885 108.535 141.160 ;
        RECT 105.610 140.605 108.980 140.885 ;
        RECT 106.080 140.295 108.980 140.605 ;
        RECT 116.450 140.870 117.050 141.170 ;
        RECT 116.450 140.570 117.350 140.870 ;
        RECT 118.250 140.570 119.150 141.470 ;
        RECT 120.350 141.170 120.650 141.470 ;
        RECT 130.425 141.305 133.100 141.860 ;
        RECT 120.350 140.870 120.950 141.170 ;
        RECT 120.050 140.570 120.950 140.870 ;
        RECT 130.765 141.135 133.100 141.305 ;
        RECT 130.765 140.585 133.425 141.135 ;
        RECT 106.080 140.040 109.415 140.295 ;
        RECT 106.535 139.700 109.415 140.040 ;
        RECT 106.535 139.465 109.840 139.700 ;
        RECT 106.980 139.095 109.840 139.465 ;
        RECT 116.450 139.370 120.950 140.570 ;
        RECT 131.100 140.405 133.425 140.585 ;
        RECT 131.100 139.860 133.745 140.405 ;
        RECT 131.425 139.670 133.745 139.860 ;
        RECT 106.980 138.885 110.255 139.095 ;
        RECT 107.415 138.480 110.255 138.885 ;
        RECT 107.415 138.295 110.660 138.480 ;
        RECT 107.840 137.865 110.660 138.295 ;
        RECT 107.840 137.700 111.055 137.865 ;
        RECT 108.255 137.350 111.055 137.700 ;
        RECT 115.170 137.780 115.730 139.170 ;
        RECT 116.750 138.770 120.650 139.370 ;
        RECT 131.425 139.135 134.050 139.670 ;
        RECT 131.745 138.930 134.050 139.135 ;
        RECT 117.350 138.470 120.050 138.770 ;
        RECT 117.650 138.170 120.050 138.470 ;
        RECT 131.745 138.405 134.350 138.930 ;
        RECT 132.050 138.190 134.350 138.405 ;
        RECT 115.170 137.350 115.620 137.780 ;
        RECT 132.050 137.670 134.635 138.190 ;
        RECT 132.350 137.530 134.635 137.670 ;
        RECT 108.255 137.095 115.620 137.350 ;
        RECT 108.660 136.900 115.620 137.095 ;
        RECT 128.900 137.445 134.635 137.530 ;
        RECT 128.900 137.080 134.915 137.445 ;
        RECT 108.660 136.605 111.440 136.900 ;
        RECT 108.660 136.480 111.810 136.605 ;
        RECT 109.055 135.970 111.810 136.480 ;
        RECT 124.470 136.300 126.870 136.600 ;
        RECT 124.470 136.000 127.170 136.300 ;
        RECT 109.055 135.865 112.170 135.970 ;
        RECT 109.440 135.325 112.170 135.865 ;
        RECT 123.870 135.400 127.770 136.000 ;
        RECT 128.900 135.530 129.350 137.080 ;
        RECT 132.350 136.930 134.915 137.080 ;
        RECT 132.635 136.695 134.915 136.930 ;
        RECT 132.635 136.190 135.185 136.695 ;
        RECT 132.915 135.940 135.185 136.190 ;
        RECT 132.915 135.445 135.445 135.940 ;
        RECT 109.440 135.240 112.520 135.325 ;
        RECT 109.810 134.675 112.520 135.240 ;
        RECT 109.810 134.605 112.860 134.675 ;
        RECT 110.170 134.020 112.860 134.605 ;
        RECT 123.570 134.200 128.070 135.400 ;
        RECT 133.185 135.185 135.445 135.445 ;
        RECT 133.185 134.695 135.695 135.185 ;
        RECT 110.170 133.970 113.185 134.020 ;
        RECT 110.520 133.355 113.185 133.970 ;
        RECT 123.570 133.900 124.470 134.200 ;
        RECT 123.570 133.600 124.170 133.900 ;
        RECT 110.520 133.325 113.500 133.355 ;
        RECT 35.075 132.620 37.695 132.675 ;
        RECT 12.490 132.135 14.710 132.430 ;
        RECT 25.360 132.170 37.695 132.620 ;
        RECT 12.275 131.665 14.710 132.135 ;
        RECT 35.075 132.020 37.695 132.170 ;
        RECT 12.275 131.365 14.490 131.665 ;
        RECT 12.075 131.360 14.490 131.365 ;
        RECT 12.075 130.910 21.250 131.360 ;
        RECT 34.780 131.355 37.380 132.020 ;
        RECT 34.780 131.340 37.075 131.355 ;
        RECT 12.075 130.900 14.490 130.910 ;
        RECT 12.075 130.590 14.275 130.900 ;
        RECT 11.880 130.135 14.275 130.590 ;
        RECT 11.880 129.815 14.075 130.135 ;
        RECT 11.695 129.365 14.075 129.815 ;
        RECT 11.695 129.040 13.880 129.365 ;
        RECT 20.800 129.360 21.250 130.910 ;
        RECT 34.500 130.690 37.075 131.340 ;
        RECT 57.540 130.730 64.170 132.940 ;
        RECT 34.500 130.660 36.780 130.690 ;
        RECT 23.280 130.130 25.680 130.430 ;
        RECT 22.980 129.830 25.680 130.130 ;
        RECT 34.230 130.020 36.780 130.660 ;
        RECT 34.230 129.970 36.500 130.020 ;
        RECT 22.380 129.230 26.280 129.830 ;
        RECT 33.975 129.340 36.500 129.970 ;
        RECT 33.975 129.280 36.230 129.340 ;
        RECT 11.525 128.590 13.880 129.040 ;
        RECT 11.525 128.260 13.695 128.590 ;
        RECT 11.360 127.815 13.695 128.260 ;
        RECT 22.080 128.030 26.580 129.230 ;
        RECT 33.730 128.660 36.230 129.280 ;
        RECT 33.730 128.585 35.975 128.660 ;
        RECT 11.360 127.480 13.525 127.815 ;
        RECT 11.205 127.040 13.525 127.480 ;
        RECT 22.080 127.730 22.980 128.030 ;
        RECT 22.080 127.430 22.680 127.730 ;
        RECT 22.380 127.130 22.680 127.430 ;
        RECT 23.880 127.130 24.780 128.030 ;
        RECT 25.680 127.730 26.580 128.030 ;
        RECT 33.500 127.970 35.975 128.585 ;
        RECT 57.540 128.520 61.960 130.730 ;
        RECT 33.500 127.885 35.730 127.970 ;
        RECT 25.980 127.430 26.580 127.730 ;
        RECT 25.980 127.130 26.280 127.430 ;
        RECT 33.280 127.280 35.730 127.885 ;
        RECT 33.280 127.185 35.500 127.280 ;
        RECT 11.205 126.695 13.360 127.040 ;
        RECT 11.060 126.260 13.360 126.695 ;
        RECT 22.380 126.830 22.980 127.130 ;
        RECT 23.580 126.830 25.080 127.130 ;
        RECT 25.680 126.830 26.280 127.130 ;
        RECT 22.380 126.530 24.180 126.830 ;
        RECT 24.480 126.530 25.980 126.830 ;
        RECT 11.060 125.910 13.205 126.260 ;
        RECT 22.980 126.230 23.880 126.530 ;
        RECT 24.780 126.230 25.980 126.530 ;
        RECT 33.070 126.585 35.500 127.185 ;
        RECT 33.070 126.480 35.280 126.585 ;
        RECT 10.925 125.480 13.205 125.910 ;
        RECT 23.280 125.630 25.380 126.230 ;
        RECT 32.875 125.885 35.280 126.480 ;
        RECT 59.750 126.310 61.960 128.520 ;
        RECT 70.800 126.310 77.430 132.940 ;
        RECT 84.060 130.730 90.690 132.940 ;
        RECT 110.860 132.690 113.500 133.325 ;
        RECT 123.870 133.300 124.170 133.600 ;
        RECT 125.370 133.300 126.270 134.200 ;
        RECT 127.170 133.900 128.070 134.200 ;
        RECT 133.445 134.430 135.695 134.695 ;
        RECT 133.445 133.940 135.940 134.430 ;
        RECT 127.470 133.600 128.070 133.900 ;
        RECT 133.695 133.665 135.940 133.940 ;
        RECT 127.470 133.300 127.770 133.600 ;
        RECT 123.870 133.000 124.470 133.300 ;
        RECT 125.070 133.000 126.570 133.300 ;
        RECT 127.170 133.000 127.770 133.300 ;
        RECT 133.695 133.185 136.170 133.665 ;
        RECT 124.170 132.700 125.670 133.000 ;
        RECT 125.970 132.700 127.770 133.000 ;
        RECT 133.940 132.900 136.170 133.185 ;
        RECT 110.860 132.675 113.805 132.690 ;
        RECT 111.185 132.020 113.805 132.675 ;
        RECT 124.170 132.400 125.370 132.700 ;
        RECT 126.270 132.400 127.170 132.700 ;
        RECT 133.940 132.430 136.390 132.900 ;
        RECT 111.500 131.355 114.100 132.020 ;
        RECT 124.770 131.800 126.870 132.400 ;
        RECT 134.170 132.135 136.390 132.430 ;
        RECT 122.970 131.500 123.870 131.800 ;
        RECT 124.770 131.500 125.070 131.800 ;
        RECT 125.370 131.500 125.670 131.800 ;
        RECT 125.970 131.500 126.270 131.800 ;
        RECT 126.570 131.500 126.870 131.800 ;
        RECT 127.770 131.500 128.670 131.800 ;
        RECT 134.170 131.665 136.605 132.135 ;
        RECT 86.270 128.520 90.690 130.730 ;
        RECT 111.805 131.340 114.100 131.355 ;
        RECT 111.805 130.690 114.380 131.340 ;
        RECT 122.670 130.900 124.170 131.500 ;
        RECT 127.470 130.900 128.970 131.500 ;
        RECT 134.390 131.365 136.605 131.665 ;
        RECT 134.390 130.900 136.805 131.365 ;
        RECT 112.100 130.660 114.380 130.690 ;
        RECT 112.100 130.020 114.650 130.660 ;
        RECT 122.970 130.600 124.770 130.900 ;
        RECT 126.870 130.600 128.670 130.900 ;
        RECT 123.870 130.300 125.070 130.600 ;
        RECT 126.570 130.300 127.770 130.600 ;
        RECT 134.605 130.590 136.805 130.900 ;
        RECT 112.380 129.970 114.650 130.020 ;
        RECT 124.470 130.000 125.670 130.300 ;
        RECT 125.970 130.000 127.170 130.300 ;
        RECT 134.605 130.135 137.000 130.590 ;
        RECT 112.380 129.340 114.905 129.970 ;
        RECT 125.070 129.400 126.570 130.000 ;
        RECT 134.805 129.815 137.000 130.135 ;
        RECT 112.650 129.280 114.905 129.340 ;
        RECT 112.650 128.660 115.150 129.280 ;
        RECT 124.470 129.100 125.670 129.400 ;
        RECT 125.970 129.100 127.170 129.400 ;
        RECT 134.805 129.365 137.185 129.815 ;
        RECT 112.905 128.585 115.150 128.660 ;
        RECT 122.670 128.800 125.070 129.100 ;
        RECT 126.570 128.800 128.670 129.100 ;
        RECT 135.000 129.040 137.185 129.365 ;
        RECT 86.270 126.310 88.480 128.520 ;
        RECT 112.905 127.970 115.380 128.585 ;
        RECT 113.150 127.885 115.380 127.970 ;
        RECT 122.670 128.500 124.470 128.800 ;
        RECT 127.170 128.500 128.970 128.800 ;
        RECT 135.000 128.590 137.355 129.040 ;
        RECT 122.670 128.200 123.870 128.500 ;
        RECT 127.770 128.200 128.970 128.500 ;
        RECT 122.670 127.900 123.570 128.200 ;
        RECT 128.070 127.900 128.970 128.200 ;
        RECT 135.185 128.260 137.355 128.590 ;
        RECT 113.150 127.280 115.600 127.885 ;
        RECT 122.970 127.600 123.270 127.900 ;
        RECT 124.770 127.600 125.070 127.900 ;
        RECT 125.370 127.600 125.670 127.900 ;
        RECT 125.970 127.600 126.270 127.900 ;
        RECT 126.570 127.600 126.870 127.900 ;
        RECT 128.370 127.600 128.670 127.900 ;
        RECT 135.185 127.815 137.520 128.260 ;
        RECT 113.380 127.185 115.600 127.280 ;
        RECT 113.380 126.585 115.810 127.185 ;
        RECT 124.770 127.000 126.870 127.600 ;
        RECT 135.355 127.480 137.520 127.815 ;
        RECT 135.355 127.040 137.675 127.480 ;
        RECT 32.875 125.770 35.070 125.885 ;
        RECT 10.925 125.125 13.060 125.480 ;
        RECT 21.480 125.330 22.380 125.630 ;
        RECT 23.280 125.330 23.580 125.630 ;
        RECT 23.880 125.330 24.180 125.630 ;
        RECT 24.480 125.330 24.780 125.630 ;
        RECT 25.080 125.330 25.380 125.630 ;
        RECT 26.280 125.330 27.180 125.630 ;
        RECT 10.800 124.695 13.060 125.125 ;
        RECT 21.180 124.730 22.680 125.330 ;
        RECT 25.980 124.730 27.480 125.330 ;
        RECT 32.690 125.185 35.070 125.770 ;
        RECT 32.690 125.055 34.875 125.185 ;
        RECT 10.800 124.340 12.925 124.695 ;
        RECT 21.480 124.430 23.280 124.730 ;
        RECT 25.380 124.430 27.180 124.730 ;
        RECT 32.520 124.480 34.875 125.055 ;
        RECT 10.685 123.910 12.925 124.340 ;
        RECT 22.380 124.130 23.580 124.430 ;
        RECT 25.080 124.130 26.280 124.430 ;
        RECT 32.520 124.340 34.690 124.480 ;
        RECT 10.685 123.550 12.800 123.910 ;
        RECT 22.980 123.830 24.180 124.130 ;
        RECT 24.480 123.830 25.680 124.130 ;
        RECT 10.580 123.125 12.800 123.550 ;
        RECT 23.580 123.230 25.080 123.830 ;
        RECT 32.360 123.770 34.690 124.340 ;
        RECT 59.750 124.100 64.170 126.310 ;
        RECT 68.590 124.100 79.640 126.310 ;
        RECT 84.060 124.100 88.480 126.310 ;
        RECT 113.600 126.480 115.810 126.585 ;
        RECT 124.170 126.700 125.370 127.000 ;
        RECT 126.270 126.700 127.170 127.000 ;
        RECT 113.600 125.885 116.005 126.480 ;
        RECT 124.170 126.400 125.670 126.700 ;
        RECT 125.970 126.400 127.770 126.700 ;
        RECT 113.810 125.770 116.005 125.885 ;
        RECT 123.870 126.100 124.470 126.400 ;
        RECT 125.070 126.100 126.570 126.400 ;
        RECT 127.170 126.100 127.770 126.400 ;
        RECT 135.520 126.695 137.675 127.040 ;
        RECT 135.520 126.260 137.820 126.695 ;
        RECT 123.870 125.800 124.170 126.100 ;
        RECT 113.810 125.185 116.190 125.770 ;
        RECT 114.005 125.055 116.190 125.185 ;
        RECT 123.570 125.500 124.170 125.800 ;
        RECT 123.570 125.200 124.470 125.500 ;
        RECT 125.370 125.200 126.270 126.100 ;
        RECT 127.470 125.800 127.770 126.100 ;
        RECT 135.675 125.910 137.820 126.260 ;
        RECT 127.470 125.500 128.070 125.800 ;
        RECT 127.170 125.200 128.070 125.500 ;
        RECT 135.675 125.480 137.955 125.910 ;
        RECT 114.005 124.480 116.360 125.055 ;
        RECT 114.190 124.340 116.360 124.480 ;
        RECT 32.360 123.620 34.520 123.770 ;
        RECT 10.580 122.760 12.685 123.125 ;
        RECT 22.980 122.930 24.180 123.230 ;
        RECT 24.480 122.930 25.680 123.230 ;
        RECT 32.215 123.055 34.520 123.620 ;
        RECT 10.485 122.340 12.685 122.760 ;
        RECT 21.480 122.630 23.580 122.930 ;
        RECT 25.080 122.630 27.480 122.930 ;
        RECT 32.215 122.900 34.360 123.055 ;
        RECT 10.485 121.965 12.580 122.340 ;
        RECT 10.400 121.550 12.580 121.965 ;
        RECT 21.180 122.330 22.980 122.630 ;
        RECT 25.680 122.330 27.480 122.630 ;
        RECT 21.180 122.030 22.380 122.330 ;
        RECT 26.280 122.030 27.480 122.330 ;
        RECT 32.080 122.340 34.360 122.900 ;
        RECT 32.080 122.180 34.215 122.340 ;
        RECT 21.180 121.730 22.080 122.030 ;
        RECT 26.580 121.730 27.480 122.030 ;
        RECT 10.400 121.175 12.485 121.550 ;
        RECT 21.480 121.430 21.780 121.730 ;
        RECT 23.280 121.430 23.580 121.730 ;
        RECT 23.880 121.430 24.180 121.730 ;
        RECT 24.480 121.430 24.780 121.730 ;
        RECT 25.080 121.430 25.380 121.730 ;
        RECT 26.880 121.430 27.180 121.730 ;
        RECT 31.960 121.620 34.215 122.180 ;
        RECT 59.750 121.890 73.010 124.100 ;
        RECT 75.220 121.890 86.270 124.100 ;
        RECT 114.190 123.770 116.520 124.340 ;
        RECT 123.570 124.000 128.070 125.200 ;
        RECT 135.820 125.125 137.955 125.480 ;
        RECT 135.820 124.695 138.080 125.125 ;
        RECT 135.955 124.340 138.080 124.695 ;
        RECT 114.360 123.620 116.520 123.770 ;
        RECT 114.360 123.055 116.665 123.620 ;
        RECT 123.870 123.400 127.770 124.000 ;
        RECT 135.955 123.910 138.195 124.340 ;
        RECT 114.520 122.900 116.665 123.055 ;
        RECT 124.470 123.100 127.170 123.400 ;
        RECT 114.520 122.340 116.800 122.900 ;
        RECT 124.470 122.800 126.870 123.100 ;
        RECT 128.790 122.410 129.350 123.800 ;
        RECT 136.080 123.550 138.195 123.910 ;
        RECT 136.080 123.125 138.300 123.550 ;
        RECT 31.960 121.455 34.080 121.620 ;
        RECT 10.325 120.760 12.485 121.175 ;
        RECT 23.280 120.830 25.380 121.430 ;
        RECT 31.850 120.900 34.080 121.455 ;
        RECT 10.325 120.380 12.400 120.760 ;
        RECT 22.980 120.530 23.880 120.830 ;
        RECT 24.780 120.530 25.980 120.830 ;
        RECT 31.850 120.725 33.960 120.900 ;
        RECT 10.265 119.965 12.400 120.380 ;
        RECT 22.380 120.230 24.180 120.530 ;
        RECT 24.480 120.230 25.980 120.530 ;
        RECT 10.265 119.585 12.325 119.965 ;
        RECT 22.380 119.930 22.980 120.230 ;
        RECT 23.580 119.930 25.080 120.230 ;
        RECT 25.680 119.930 26.280 120.230 ;
        RECT 31.755 120.180 33.960 120.725 ;
        RECT 31.755 120.000 33.850 120.180 ;
        RECT 22.380 119.630 22.680 119.930 ;
        RECT 10.210 119.175 12.325 119.585 ;
        RECT 22.080 119.330 22.680 119.630 ;
        RECT 10.210 118.790 12.265 119.175 ;
        RECT 10.165 118.380 12.265 118.790 ;
        RECT 22.080 119.030 22.980 119.330 ;
        RECT 23.880 119.030 24.780 119.930 ;
        RECT 25.980 119.630 26.280 119.930 ;
        RECT 25.980 119.330 26.580 119.630 ;
        RECT 25.680 119.030 26.580 119.330 ;
        RECT 31.675 119.455 33.850 120.000 ;
        RECT 64.170 119.680 70.800 121.890 ;
        RECT 77.430 119.680 86.270 121.890 ;
        RECT 114.665 122.180 116.800 122.340 ;
        RECT 114.665 121.980 116.920 122.180 ;
        RECT 128.900 121.980 129.350 122.410 ;
        RECT 136.195 122.760 138.300 123.125 ;
        RECT 136.195 122.340 138.395 122.760 ;
        RECT 114.665 121.620 129.350 121.980 ;
        RECT 114.800 121.530 129.350 121.620 ;
        RECT 136.300 121.965 138.395 122.340 ;
        RECT 136.300 121.550 138.480 121.965 ;
        RECT 114.800 121.145 117.175 121.530 ;
        RECT 136.395 121.175 138.480 121.550 ;
        RECT 114.800 120.900 117.030 121.145 ;
        RECT 114.920 120.725 117.030 120.900 ;
        RECT 136.395 120.760 138.555 121.175 ;
        RECT 114.920 120.180 117.125 120.725 ;
        RECT 136.480 120.610 138.555 120.760 ;
        RECT 115.030 120.000 117.125 120.180 ;
        RECT 126.210 120.380 138.555 120.610 ;
        RECT 126.210 120.160 138.615 120.380 ;
        RECT 31.675 119.270 33.755 119.455 ;
        RECT 10.165 117.995 12.210 118.380 ;
        RECT 10.130 117.585 12.210 117.995 ;
        RECT 22.080 117.830 26.580 119.030 ;
        RECT 31.600 118.725 33.755 119.270 ;
        RECT 31.600 118.535 33.675 118.725 ;
        RECT 31.545 118.000 33.675 118.535 ;
        RECT 10.130 117.200 12.165 117.585 ;
        RECT 10.105 116.790 12.165 117.200 ;
        RECT 10.105 116.405 12.130 116.790 ;
        RECT 10.090 115.995 12.130 116.405 ;
        RECT 20.800 116.240 21.360 117.630 ;
        RECT 22.380 117.230 26.280 117.830 ;
        RECT 31.545 117.805 33.600 118.000 ;
        RECT 31.500 117.270 33.600 117.805 ;
        RECT 22.980 116.930 25.680 117.230 ;
        RECT 31.500 117.075 33.545 117.270 ;
        RECT 23.280 116.630 25.680 116.930 ;
        RECT 31.470 116.535 33.545 117.075 ;
        RECT 31.470 116.340 33.500 116.535 ;
        RECT 10.090 115.610 12.105 115.995 ;
        RECT 10.080 115.200 12.105 115.610 ;
        RECT 20.800 115.810 21.250 116.240 ;
        RECT 31.450 115.810 33.500 116.340 ;
        RECT 20.800 115.805 33.500 115.810 ;
        RECT 20.800 115.360 33.470 115.805 ;
        RECT 10.080 114.860 12.090 115.200 ;
        RECT 31.440 115.075 33.470 115.360 ;
        RECT 66.380 115.260 81.850 119.680 ;
        RECT 115.030 119.455 117.205 120.000 ;
        RECT 115.125 119.270 117.205 119.455 ;
        RECT 115.125 118.725 117.280 119.270 ;
        RECT 115.205 118.535 117.280 118.725 ;
        RECT 126.210 118.610 126.660 120.160 ;
        RECT 136.480 119.965 138.615 120.160 ;
        RECT 128.690 119.380 131.090 119.680 ;
        RECT 128.390 119.080 131.090 119.380 ;
        RECT 136.555 119.585 138.615 119.965 ;
        RECT 136.555 119.175 138.670 119.585 ;
        RECT 115.205 118.000 117.335 118.535 ;
        RECT 127.790 118.480 131.690 119.080 ;
        RECT 136.615 118.790 138.670 119.175 ;
        RECT 115.280 117.805 117.335 118.000 ;
        RECT 115.280 117.270 117.380 117.805 ;
        RECT 115.335 117.075 117.380 117.270 ;
        RECT 127.490 117.280 131.990 118.480 ;
        RECT 136.615 118.380 138.715 118.790 ;
        RECT 136.670 117.995 138.715 118.380 ;
        RECT 136.670 117.585 138.750 117.995 ;
        RECT 115.335 116.535 117.410 117.075 ;
        RECT 127.490 116.980 128.390 117.280 ;
        RECT 127.490 116.680 128.090 116.980 ;
        RECT 115.380 116.340 117.410 116.535 ;
        RECT 127.790 116.380 128.090 116.680 ;
        RECT 129.290 116.380 130.190 117.280 ;
        RECT 131.090 116.980 131.990 117.280 ;
        RECT 131.390 116.680 131.990 116.980 ;
        RECT 136.715 117.200 138.750 117.585 ;
        RECT 136.715 116.790 138.775 117.200 ;
        RECT 131.390 116.380 131.690 116.680 ;
        RECT 115.380 115.805 117.430 116.340 ;
        RECT 115.410 115.610 117.430 115.805 ;
        RECT 127.790 116.080 128.390 116.380 ;
        RECT 128.990 116.080 130.490 116.380 ;
        RECT 131.090 116.080 131.690 116.380 ;
        RECT 136.750 116.405 138.775 116.790 ;
        RECT 127.790 115.780 129.590 116.080 ;
        RECT 129.890 115.780 131.390 116.080 ;
        RECT 136.750 115.995 138.790 116.405 ;
        RECT 7.520 114.410 9.020 114.460 ;
        RECT 10.080 114.410 17.250 114.860 ;
        RECT 7.520 114.020 12.090 114.410 ;
        RECT 7.520 113.225 12.105 114.020 ;
        RECT 7.520 112.910 12.130 113.225 ;
        RECT 7.520 112.860 9.020 112.910 ;
        RECT 10.090 112.815 12.130 112.910 ;
        RECT 16.800 112.860 17.250 114.410 ;
        RECT 31.440 114.145 33.450 115.075 ;
        RECT 19.280 113.630 21.680 113.930 ;
        RECT 18.980 113.330 21.680 113.630 ;
        RECT 31.440 113.615 33.470 114.145 ;
        RECT 31.450 113.415 33.470 113.615 ;
        RECT 10.105 112.430 12.130 112.815 ;
        RECT 18.380 112.730 22.280 113.330 ;
        RECT 31.450 112.880 33.500 113.415 ;
        RECT 53.120 113.050 59.750 115.260 ;
        RECT 66.380 113.050 68.590 115.260 ;
        RECT 70.800 113.050 73.010 115.260 ;
        RECT 75.220 113.050 77.430 115.260 ;
        RECT 79.640 113.050 81.850 115.260 ;
        RECT 88.480 113.050 95.110 115.260 ;
        RECT 115.410 115.075 117.440 115.610 ;
        RECT 128.390 115.480 129.290 115.780 ;
        RECT 130.190 115.480 131.390 115.780 ;
        RECT 136.775 115.610 138.790 115.995 ;
        RECT 115.430 114.145 117.440 115.075 ;
        RECT 128.690 114.880 130.790 115.480 ;
        RECT 136.775 115.200 138.800 115.610 ;
        RECT 126.890 114.580 127.790 114.880 ;
        RECT 128.690 114.580 128.990 114.880 ;
        RECT 129.290 114.580 129.590 114.880 ;
        RECT 129.890 114.580 130.190 114.880 ;
        RECT 130.490 114.580 130.790 114.880 ;
        RECT 131.690 114.580 132.590 114.880 ;
        RECT 115.410 113.610 117.440 114.145 ;
        RECT 126.590 113.980 128.090 114.580 ;
        RECT 131.390 113.980 132.890 114.580 ;
        RECT 136.790 114.020 138.800 115.200 ;
        RECT 126.890 113.680 128.690 113.980 ;
        RECT 130.790 113.680 132.590 113.980 ;
        RECT 115.410 113.415 117.430 113.610 ;
        RECT 10.105 112.020 12.165 112.430 ;
        RECT 10.130 111.635 12.165 112.020 ;
        RECT 10.130 111.225 12.210 111.635 ;
        RECT 10.165 110.840 12.210 111.225 ;
        RECT 18.080 111.530 22.580 112.730 ;
        RECT 31.470 112.685 33.500 112.880 ;
        RECT 31.470 112.145 33.545 112.685 ;
        RECT 18.080 111.230 18.980 111.530 ;
        RECT 18.080 110.930 18.680 111.230 ;
        RECT 10.165 110.430 12.265 110.840 ;
        RECT 10.210 110.045 12.265 110.430 ;
        RECT 18.380 110.630 18.680 110.930 ;
        RECT 19.880 110.630 20.780 111.530 ;
        RECT 21.680 111.230 22.580 111.530 ;
        RECT 31.500 111.950 33.545 112.145 ;
        RECT 31.500 111.415 33.600 111.950 ;
        RECT 21.980 110.930 22.580 111.230 ;
        RECT 31.545 111.220 33.600 111.415 ;
        RECT 21.980 110.630 22.280 110.930 ;
        RECT 31.545 110.685 33.675 111.220 ;
        RECT 18.380 110.330 18.980 110.630 ;
        RECT 19.580 110.330 21.080 110.630 ;
        RECT 21.680 110.330 22.280 110.630 ;
        RECT 31.600 110.495 33.675 110.685 ;
        RECT 10.210 109.635 12.325 110.045 ;
        RECT 18.380 110.030 20.180 110.330 ;
        RECT 20.480 110.030 21.980 110.330 ;
        RECT 18.980 109.730 19.880 110.030 ;
        RECT 20.780 109.730 21.980 110.030 ;
        RECT 31.600 109.950 33.755 110.495 ;
        RECT 31.675 109.765 33.755 109.950 ;
        RECT 10.265 109.255 12.325 109.635 ;
        RECT 10.265 108.840 12.400 109.255 ;
        RECT 19.280 109.130 21.380 109.730 ;
        RECT 31.675 109.220 33.850 109.765 ;
        RECT 10.325 108.460 12.400 108.840 ;
        RECT 17.480 108.830 18.380 109.130 ;
        RECT 19.280 108.830 19.580 109.130 ;
        RECT 19.880 108.830 20.180 109.130 ;
        RECT 20.480 108.830 20.780 109.130 ;
        RECT 21.080 108.830 21.380 109.130 ;
        RECT 22.280 108.830 23.180 109.130 ;
        RECT 31.755 109.040 33.850 109.220 ;
        RECT 10.325 108.045 12.485 108.460 ;
        RECT 17.180 108.230 18.680 108.830 ;
        RECT 21.980 108.230 23.480 108.830 ;
        RECT 31.755 108.495 33.960 109.040 ;
        RECT 50.910 108.630 61.960 113.050 ;
        RECT 86.270 108.630 97.320 113.050 ;
        RECT 115.380 112.880 117.430 113.415 ;
        RECT 127.790 113.380 128.990 113.680 ;
        RECT 130.490 113.380 131.690 113.680 ;
        RECT 136.775 113.610 138.800 114.020 ;
        RECT 128.390 113.080 129.590 113.380 ;
        RECT 129.890 113.080 131.090 113.380 ;
        RECT 136.775 113.225 138.790 113.610 ;
        RECT 115.380 112.685 117.410 112.880 ;
        RECT 115.335 112.145 117.410 112.685 ;
        RECT 128.990 112.480 130.490 113.080 ;
        RECT 136.750 112.815 138.790 113.225 ;
        RECT 128.390 112.180 129.590 112.480 ;
        RECT 129.890 112.180 131.090 112.480 ;
        RECT 136.750 112.430 138.775 112.815 ;
        RECT 115.335 111.950 117.380 112.145 ;
        RECT 115.280 111.415 117.380 111.950 ;
        RECT 126.890 111.880 128.990 112.180 ;
        RECT 130.490 111.880 132.890 112.180 ;
        RECT 126.590 111.580 128.390 111.880 ;
        RECT 131.090 111.580 132.890 111.880 ;
        RECT 136.715 112.020 138.775 112.430 ;
        RECT 136.715 111.635 138.750 112.020 ;
        RECT 115.280 111.220 117.335 111.415 ;
        RECT 115.205 110.685 117.335 111.220 ;
        RECT 126.590 111.280 127.790 111.580 ;
        RECT 131.690 111.280 132.890 111.580 ;
        RECT 126.590 110.980 127.490 111.280 ;
        RECT 131.990 110.980 132.890 111.280 ;
        RECT 136.670 111.225 138.750 111.635 ;
        RECT 115.205 110.495 117.280 110.685 ;
        RECT 126.890 110.680 127.190 110.980 ;
        RECT 128.690 110.680 128.990 110.980 ;
        RECT 129.290 110.680 129.590 110.980 ;
        RECT 129.890 110.680 130.190 110.980 ;
        RECT 130.490 110.680 130.790 110.980 ;
        RECT 132.290 110.680 132.590 110.980 ;
        RECT 136.670 110.840 138.715 111.225 ;
        RECT 115.125 109.950 117.280 110.495 ;
        RECT 128.690 110.080 130.790 110.680 ;
        RECT 136.615 110.430 138.715 110.840 ;
        RECT 115.125 109.765 117.205 109.950 ;
        RECT 128.390 109.780 129.290 110.080 ;
        RECT 130.190 109.780 131.390 110.080 ;
        RECT 136.615 110.045 138.670 110.430 ;
        RECT 115.030 109.220 117.205 109.765 ;
        RECT 127.790 109.480 129.590 109.780 ;
        RECT 129.890 109.480 131.390 109.780 ;
        RECT 136.555 109.635 138.670 110.045 ;
        RECT 115.030 109.040 117.125 109.220 ;
        RECT 31.850 108.320 33.960 108.495 ;
        RECT 10.400 107.670 12.485 108.045 ;
        RECT 17.480 107.930 19.280 108.230 ;
        RECT 21.380 107.930 23.180 108.230 ;
        RECT 10.400 107.255 12.580 107.670 ;
        RECT 18.380 107.630 19.580 107.930 ;
        RECT 21.080 107.630 22.280 107.930 ;
        RECT 31.850 107.765 34.080 108.320 ;
        RECT 18.980 107.330 20.180 107.630 ;
        RECT 20.480 107.330 21.680 107.630 ;
        RECT 31.960 107.600 34.080 107.765 ;
        RECT 10.485 106.880 12.580 107.255 ;
        RECT 10.485 106.460 12.685 106.880 ;
        RECT 19.580 106.730 21.080 107.330 ;
        RECT 31.960 107.040 34.215 107.600 ;
        RECT 32.080 106.880 34.215 107.040 ;
        RECT 10.580 106.095 12.685 106.460 ;
        RECT 18.980 106.430 20.180 106.730 ;
        RECT 20.480 106.430 21.680 106.730 ;
        RECT 17.480 106.130 19.580 106.430 ;
        RECT 21.080 106.130 23.480 106.430 ;
        RECT 32.080 106.320 34.360 106.880 ;
        RECT 53.120 106.420 66.380 108.630 ;
        RECT 81.850 106.420 95.110 108.630 ;
        RECT 114.920 108.495 117.125 109.040 ;
        RECT 127.790 109.180 128.390 109.480 ;
        RECT 128.990 109.180 130.490 109.480 ;
        RECT 131.090 109.180 131.690 109.480 ;
        RECT 136.555 109.255 138.615 109.635 ;
        RECT 127.790 108.880 128.090 109.180 ;
        RECT 127.490 108.580 128.090 108.880 ;
        RECT 114.920 108.320 117.030 108.495 ;
        RECT 114.800 107.765 117.030 108.320 ;
        RECT 127.490 108.280 128.390 108.580 ;
        RECT 129.290 108.280 130.190 109.180 ;
        RECT 131.390 108.880 131.690 109.180 ;
        RECT 131.390 108.580 131.990 108.880 ;
        RECT 131.090 108.280 131.990 108.580 ;
        RECT 136.480 108.840 138.615 109.255 ;
        RECT 136.480 108.460 138.555 108.840 ;
        RECT 114.800 107.600 116.920 107.765 ;
        RECT 114.665 107.040 116.920 107.600 ;
        RECT 127.490 107.080 131.990 108.280 ;
        RECT 136.395 108.045 138.555 108.460 ;
        RECT 136.395 107.670 138.480 108.045 ;
        RECT 136.300 107.255 138.480 107.670 ;
        RECT 114.665 106.880 116.800 107.040 ;
        RECT 10.580 105.670 12.800 106.095 ;
        RECT 10.685 105.310 12.800 105.670 ;
        RECT 17.180 105.830 18.980 106.130 ;
        RECT 21.680 105.830 23.480 106.130 ;
        RECT 17.180 105.530 18.380 105.830 ;
        RECT 22.280 105.530 23.480 105.830 ;
        RECT 32.215 106.165 34.360 106.320 ;
        RECT 32.215 105.600 34.520 106.165 ;
        RECT 10.685 104.880 12.925 105.310 ;
        RECT 17.180 105.230 18.080 105.530 ;
        RECT 22.580 105.230 23.480 105.530 ;
        RECT 32.360 105.450 34.520 105.600 ;
        RECT 17.480 104.930 17.780 105.230 ;
        RECT 19.280 104.930 19.580 105.230 ;
        RECT 19.880 104.930 20.180 105.230 ;
        RECT 20.480 104.930 20.780 105.230 ;
        RECT 21.080 104.930 21.380 105.230 ;
        RECT 22.880 104.930 23.180 105.230 ;
        RECT 10.800 104.525 12.925 104.880 ;
        RECT 10.800 104.095 13.060 104.525 ;
        RECT 19.280 104.330 21.380 104.930 ;
        RECT 32.360 104.880 34.690 105.450 ;
        RECT 32.520 104.740 34.690 104.880 ;
        RECT 10.925 103.740 13.060 104.095 ;
        RECT 18.980 104.030 19.880 104.330 ;
        RECT 20.780 104.030 21.980 104.330 ;
        RECT 32.520 104.165 34.875 104.740 ;
        RECT 59.750 104.210 68.590 106.420 ;
        RECT 79.640 104.210 88.480 106.420 ;
        RECT 114.520 106.320 116.800 106.880 ;
        RECT 114.520 106.165 116.665 106.320 ;
        RECT 114.360 105.600 116.665 106.165 ;
        RECT 114.360 105.450 116.520 105.600 ;
        RECT 114.190 105.060 116.520 105.450 ;
        RECT 126.210 105.490 126.770 106.880 ;
        RECT 127.790 106.480 131.690 107.080 ;
        RECT 136.300 106.880 138.395 107.255 ;
        RECT 128.390 106.180 131.090 106.480 ;
        RECT 128.690 105.880 131.090 106.180 ;
        RECT 136.195 106.460 138.395 106.880 ;
        RECT 136.195 106.095 138.300 106.460 ;
        RECT 136.080 105.670 138.300 106.095 ;
        RECT 126.210 105.065 126.660 105.490 ;
        RECT 136.080 105.310 138.195 105.670 ;
        RECT 125.555 105.060 129.110 105.065 ;
        RECT 114.190 104.740 129.110 105.060 ;
        RECT 114.005 104.615 129.110 104.740 ;
        RECT 114.005 104.610 126.660 104.615 ;
        RECT 10.925 103.310 13.205 103.740 ;
        RECT 11.060 102.960 13.205 103.310 ;
        RECT 18.380 103.730 20.180 104.030 ;
        RECT 20.480 103.730 21.980 104.030 ;
        RECT 32.690 104.035 34.875 104.165 ;
        RECT 18.380 103.430 18.980 103.730 ;
        RECT 19.580 103.430 21.080 103.730 ;
        RECT 21.680 103.430 22.280 103.730 ;
        RECT 32.690 103.450 35.070 104.035 ;
        RECT 18.380 103.130 18.680 103.430 ;
        RECT 11.060 102.525 13.360 102.960 ;
        RECT 11.205 102.180 13.360 102.525 ;
        RECT 18.080 102.830 18.680 103.130 ;
        RECT 18.080 102.530 18.980 102.830 ;
        RECT 19.880 102.530 20.780 103.430 ;
        RECT 21.980 103.130 22.280 103.430 ;
        RECT 32.875 103.335 35.070 103.450 ;
        RECT 21.980 102.830 22.580 103.130 ;
        RECT 21.680 102.530 22.580 102.830 ;
        RECT 32.875 102.740 35.280 103.335 ;
        RECT 11.205 101.740 13.525 102.180 ;
        RECT 11.360 101.405 13.525 101.740 ;
        RECT 11.360 100.960 13.695 101.405 ;
        RECT 18.080 101.330 22.580 102.530 ;
        RECT 33.070 102.635 35.280 102.740 ;
        RECT 33.070 102.035 35.500 102.635 ;
        RECT 33.280 101.940 35.500 102.035 ;
        RECT 64.170 102.000 73.010 104.210 ;
        RECT 75.220 102.000 84.060 104.210 ;
        RECT 114.005 104.165 116.360 104.610 ;
        RECT 114.005 104.035 116.190 104.165 ;
        RECT 113.810 103.450 116.190 104.035 ;
        RECT 113.810 103.335 116.005 103.450 ;
        RECT 113.600 102.740 116.005 103.335 ;
        RECT 128.660 102.860 129.110 104.615 ;
        RECT 135.955 104.880 138.195 105.310 ;
        RECT 135.955 104.525 138.080 104.880 ;
        RECT 135.820 104.095 138.080 104.525 ;
        RECT 135.820 103.740 137.955 104.095 ;
        RECT 135.675 103.310 137.955 103.740 ;
        RECT 135.675 102.960 137.820 103.310 ;
        RECT 113.600 102.635 115.810 102.740 ;
        RECT 113.380 102.035 115.810 102.635 ;
        RECT 124.190 102.170 126.590 102.470 ;
        RECT 128.510 102.290 129.110 102.860 ;
        RECT 135.520 102.525 137.820 102.960 ;
        RECT 33.280 101.335 35.730 101.940 ;
        RECT 11.525 100.630 13.695 100.960 ;
        RECT 11.525 100.180 13.880 100.630 ;
        RECT 11.695 99.855 13.880 100.180 ;
        RECT 11.695 99.405 14.075 99.855 ;
        RECT 11.880 99.085 14.075 99.405 ;
        RECT 16.800 99.740 17.360 101.130 ;
        RECT 18.380 100.730 22.280 101.330 ;
        RECT 33.500 101.250 35.730 101.335 ;
        RECT 18.980 100.430 21.680 100.730 ;
        RECT 33.500 100.635 35.975 101.250 ;
        RECT 19.280 100.130 21.680 100.430 ;
        RECT 33.730 100.560 35.975 100.635 ;
        RECT 33.730 99.940 36.230 100.560 ;
        RECT 33.975 99.880 36.230 99.940 ;
        RECT 16.800 99.315 17.250 99.740 ;
        RECT 33.975 99.315 36.500 99.880 ;
        RECT 16.800 99.200 36.500 99.315 ;
        RECT 11.880 98.630 14.275 99.085 ;
        RECT 16.800 98.865 36.780 99.200 ;
        RECT 16.800 98.860 17.250 98.865 ;
        RECT 12.075 98.320 14.275 98.630 ;
        RECT 34.230 98.560 36.780 98.865 ;
        RECT 34.500 98.530 36.780 98.560 ;
        RECT 12.075 98.175 14.490 98.320 ;
        RECT 12.075 97.855 29.320 98.175 ;
        RECT 34.500 97.880 37.075 98.530 ;
        RECT 12.275 97.725 29.320 97.855 ;
        RECT 12.275 97.555 14.490 97.725 ;
        RECT 12.275 97.085 14.710 97.555 ;
        RECT 12.490 96.790 14.710 97.085 ;
        RECT 24.440 96.820 26.840 97.120 ;
        RECT 12.490 96.320 14.940 96.790 ;
        RECT 24.440 96.520 27.140 96.820 ;
        RECT 12.710 96.035 14.940 96.320 ;
        RECT 12.710 95.555 15.185 96.035 ;
        RECT 23.840 95.920 27.740 96.520 ;
        RECT 28.870 96.050 29.320 97.725 ;
        RECT 34.780 97.865 37.075 97.880 ;
        RECT 34.780 97.200 37.380 97.865 ;
        RECT 68.590 97.580 79.640 102.000 ;
        RECT 113.380 101.940 115.600 102.035 ;
        RECT 113.150 101.335 115.600 101.940 ;
        RECT 124.190 101.870 126.890 102.170 ;
        RECT 113.150 101.250 115.380 101.335 ;
        RECT 123.590 101.270 127.490 101.870 ;
        RECT 128.510 101.470 129.070 102.290 ;
        RECT 135.520 102.180 137.675 102.525 ;
        RECT 135.355 101.740 137.675 102.180 ;
        RECT 135.355 101.405 137.520 101.740 ;
        RECT 112.905 100.635 115.380 101.250 ;
        RECT 112.905 100.560 115.150 100.635 ;
        RECT 112.650 99.940 115.150 100.560 ;
        RECT 123.290 100.070 127.790 101.270 ;
        RECT 135.185 100.960 137.520 101.405 ;
        RECT 135.185 100.630 137.355 100.960 ;
        RECT 112.650 99.880 114.905 99.940 ;
        RECT 112.380 99.250 114.905 99.880 ;
        RECT 123.290 99.770 124.190 100.070 ;
        RECT 123.290 99.470 123.890 99.770 ;
        RECT 112.380 99.200 114.650 99.250 ;
        RECT 112.100 98.560 114.650 99.200 ;
        RECT 123.590 99.170 123.890 99.470 ;
        RECT 125.090 99.170 125.990 100.070 ;
        RECT 126.890 99.770 127.790 100.070 ;
        RECT 135.000 100.180 137.355 100.630 ;
        RECT 135.000 99.855 137.185 100.180 ;
        RECT 127.190 99.470 127.790 99.770 ;
        RECT 127.190 99.170 127.490 99.470 ;
        RECT 123.590 98.870 124.190 99.170 ;
        RECT 124.790 98.870 126.290 99.170 ;
        RECT 126.890 98.870 127.490 99.170 ;
        RECT 134.805 99.405 137.185 99.855 ;
        RECT 134.805 99.085 137.000 99.405 ;
        RECT 123.890 98.570 125.390 98.870 ;
        RECT 125.690 98.570 127.490 98.870 ;
        RECT 134.605 98.630 137.000 99.085 ;
        RECT 112.100 98.530 114.380 98.560 ;
        RECT 111.805 97.880 114.380 98.530 ;
        RECT 123.890 98.270 125.090 98.570 ;
        RECT 125.990 98.270 126.890 98.570 ;
        RECT 134.605 98.320 136.805 98.630 ;
        RECT 111.805 97.865 114.100 97.880 ;
        RECT 35.075 96.545 37.695 97.200 ;
        RECT 35.075 96.530 38.020 96.545 ;
        RECT 12.940 95.280 15.185 95.555 ;
        RECT 12.940 94.790 15.435 95.280 ;
        RECT 13.185 94.525 15.435 94.790 ;
        RECT 23.540 94.720 28.040 95.920 ;
        RECT 35.380 95.895 38.020 96.530 ;
        RECT 35.380 95.865 38.360 95.895 ;
        RECT 35.695 95.250 38.360 95.865 ;
        RECT 64.170 95.370 73.010 97.580 ;
        RECT 75.220 95.370 84.060 97.580 ;
        RECT 111.500 97.200 114.100 97.865 ;
        RECT 124.490 97.670 126.590 98.270 ;
        RECT 134.390 97.855 136.805 98.320 ;
        RECT 122.690 97.370 122.990 97.670 ;
        RECT 124.490 97.370 124.790 97.670 ;
        RECT 125.090 97.370 125.390 97.670 ;
        RECT 125.690 97.370 125.990 97.670 ;
        RECT 126.290 97.370 126.590 97.670 ;
        RECT 128.090 97.370 128.390 97.670 ;
        RECT 134.390 97.555 136.605 97.855 ;
        RECT 111.185 96.545 113.805 97.200 ;
        RECT 110.860 96.530 113.805 96.545 ;
        RECT 122.390 97.070 123.290 97.370 ;
        RECT 127.790 97.070 128.690 97.370 ;
        RECT 122.390 96.770 123.590 97.070 ;
        RECT 127.490 96.770 128.690 97.070 ;
        RECT 134.170 97.085 136.605 97.555 ;
        RECT 134.170 96.790 136.390 97.085 ;
        RECT 110.860 95.895 113.500 96.530 ;
        RECT 122.390 96.470 124.190 96.770 ;
        RECT 126.890 96.470 128.690 96.770 ;
        RECT 122.390 96.170 124.790 96.470 ;
        RECT 126.290 96.170 128.390 96.470 ;
        RECT 133.940 96.320 136.390 96.790 ;
        RECT 110.520 95.865 113.500 95.895 ;
        RECT 124.190 95.870 125.390 96.170 ;
        RECT 125.690 95.870 126.890 96.170 ;
        RECT 133.940 96.035 136.170 96.320 ;
        RECT 35.695 95.200 38.710 95.250 ;
        RECT 13.185 94.035 15.695 94.525 ;
        RECT 23.540 94.420 24.440 94.720 ;
        RECT 23.540 94.120 24.140 94.420 ;
        RECT 13.435 93.775 15.695 94.035 ;
        RECT 23.840 93.820 24.140 94.120 ;
        RECT 25.340 93.820 26.240 94.720 ;
        RECT 27.140 94.420 28.040 94.720 ;
        RECT 36.020 94.610 38.710 95.200 ;
        RECT 36.020 94.545 39.070 94.610 ;
        RECT 27.440 94.120 28.040 94.420 ;
        RECT 27.440 93.820 27.740 94.120 ;
        RECT 36.360 93.980 39.070 94.545 ;
        RECT 36.360 93.895 39.440 93.980 ;
        RECT 13.435 93.280 15.965 93.775 ;
        RECT 23.840 93.520 24.440 93.820 ;
        RECT 25.040 93.520 26.540 93.820 ;
        RECT 27.140 93.520 27.740 93.820 ;
        RECT 13.695 93.030 15.965 93.280 ;
        RECT 24.140 93.220 25.640 93.520 ;
        RECT 25.940 93.220 27.740 93.520 ;
        RECT 36.710 93.355 39.440 93.895 ;
        RECT 36.710 93.250 39.825 93.355 ;
        RECT 13.695 92.525 16.245 93.030 ;
        RECT 24.140 92.920 25.340 93.220 ;
        RECT 26.240 92.920 27.140 93.220 ;
        RECT 13.965 92.290 16.245 92.525 ;
        RECT 24.740 92.320 26.840 92.920 ;
        RECT 37.070 92.740 39.825 93.250 ;
        RECT 53.120 93.160 68.590 95.370 ;
        RECT 79.640 93.160 97.320 95.370 ;
        RECT 110.520 95.250 113.185 95.865 ;
        RECT 124.790 95.270 126.290 95.870 ;
        RECT 133.695 95.555 136.170 96.035 ;
        RECT 133.695 95.280 135.940 95.555 ;
        RECT 110.170 95.200 113.185 95.250 ;
        RECT 110.170 94.610 112.860 95.200 ;
        RECT 124.190 94.970 125.390 95.270 ;
        RECT 125.690 94.970 126.890 95.270 ;
        RECT 123.590 94.670 124.790 94.970 ;
        RECT 126.290 94.670 127.490 94.970 ;
        RECT 133.445 94.790 135.940 95.280 ;
        RECT 109.810 94.545 112.860 94.610 ;
        RECT 109.810 93.980 112.520 94.545 ;
        RECT 122.690 94.370 124.490 94.670 ;
        RECT 126.590 94.370 128.390 94.670 ;
        RECT 133.445 94.525 135.695 94.790 ;
        RECT 109.440 93.895 112.520 93.980 ;
        RECT 109.440 93.355 112.170 93.895 ;
        RECT 122.390 93.770 123.890 94.370 ;
        RECT 127.190 93.770 128.690 94.370 ;
        RECT 133.185 94.035 135.695 94.525 ;
        RECT 133.185 93.775 135.445 94.035 ;
        RECT 122.690 93.470 123.590 93.770 ;
        RECT 124.490 93.470 124.790 93.770 ;
        RECT 125.090 93.470 125.390 93.770 ;
        RECT 125.690 93.470 125.990 93.770 ;
        RECT 126.290 93.470 126.590 93.770 ;
        RECT 127.490 93.470 128.390 93.770 ;
        RECT 37.070 92.610 40.220 92.740 ;
        RECT 13.965 91.775 16.530 92.290 ;
        RECT 22.940 92.020 23.840 92.320 ;
        RECT 24.740 92.020 25.040 92.320 ;
        RECT 25.340 92.020 25.640 92.320 ;
        RECT 25.940 92.020 26.240 92.320 ;
        RECT 26.540 92.020 26.840 92.320 ;
        RECT 27.740 92.020 28.640 92.320 ;
        RECT 37.440 92.125 40.220 92.610 ;
        RECT 14.245 91.550 16.530 91.775 ;
        RECT 14.245 91.030 16.830 91.550 ;
        RECT 22.640 91.420 24.140 92.020 ;
        RECT 27.440 91.420 28.940 92.020 ;
        RECT 37.440 91.980 40.625 92.125 ;
        RECT 37.825 91.520 40.625 91.980 ;
        RECT 22.940 91.120 24.740 91.420 ;
        RECT 26.840 91.120 28.640 91.420 ;
        RECT 37.825 91.355 41.040 91.520 ;
        RECT 14.530 90.815 16.830 91.030 ;
        RECT 23.840 90.820 25.040 91.120 ;
        RECT 26.540 90.820 27.740 91.120 ;
        RECT 38.220 90.925 41.040 91.355 ;
        RECT 50.910 90.950 64.170 93.160 ;
        RECT 84.060 90.950 97.320 93.160 ;
        RECT 109.055 93.250 112.170 93.355 ;
        RECT 109.055 92.740 111.810 93.250 ;
        RECT 124.490 92.870 126.590 93.470 ;
        RECT 132.915 93.280 135.445 93.775 ;
        RECT 132.915 93.030 135.185 93.280 ;
        RECT 108.660 92.610 111.810 92.740 ;
        RECT 108.660 92.125 111.440 92.610 ;
        RECT 123.890 92.570 125.090 92.870 ;
        RECT 125.990 92.570 126.890 92.870 ;
        RECT 123.890 92.270 125.390 92.570 ;
        RECT 125.690 92.270 127.490 92.570 ;
        RECT 132.635 92.525 135.185 93.030 ;
        RECT 132.635 92.290 134.915 92.525 ;
        RECT 108.255 91.980 111.440 92.125 ;
        RECT 108.255 91.520 111.055 91.980 ;
        RECT 123.590 91.970 124.190 92.270 ;
        RECT 124.790 91.970 126.290 92.270 ;
        RECT 126.890 91.970 127.490 92.270 ;
        RECT 123.590 91.670 123.890 91.970 ;
        RECT 14.530 90.290 17.135 90.815 ;
        RECT 24.440 90.520 25.640 90.820 ;
        RECT 25.940 90.520 27.140 90.820 ;
        RECT 38.220 90.740 41.465 90.925 ;
        RECT 14.830 90.085 17.135 90.290 ;
        RECT 14.830 89.550 17.455 90.085 ;
        RECT 25.040 89.920 26.540 90.520 ;
        RECT 38.625 90.335 41.465 90.740 ;
        RECT 38.625 90.125 41.900 90.335 ;
        RECT 24.440 89.620 25.640 89.920 ;
        RECT 25.940 89.620 27.140 89.920 ;
        RECT 39.040 89.915 41.900 90.125 ;
        RECT 38.110 89.755 41.900 89.915 ;
        RECT 15.135 89.360 17.455 89.550 ;
        RECT 15.135 88.815 17.780 89.360 ;
        RECT 15.455 88.635 17.780 88.815 ;
        RECT 22.640 89.320 25.040 89.620 ;
        RECT 26.540 89.320 28.640 89.620 ;
        RECT 38.110 89.465 42.345 89.755 ;
        RECT 22.640 89.020 24.440 89.320 ;
        RECT 27.140 89.020 28.940 89.320 ;
        RECT 22.640 88.720 23.840 89.020 ;
        RECT 27.740 88.720 28.940 89.020 ;
        RECT 15.455 88.085 18.115 88.635 ;
        RECT 22.640 88.420 23.540 88.720 ;
        RECT 28.040 88.420 28.940 88.720 ;
        RECT 22.940 88.120 23.240 88.420 ;
        RECT 24.740 88.120 25.040 88.420 ;
        RECT 25.340 88.120 25.640 88.420 ;
        RECT 25.940 88.120 26.240 88.420 ;
        RECT 26.540 88.120 26.840 88.420 ;
        RECT 28.340 88.120 28.640 88.420 ;
        RECT 15.780 87.915 18.115 88.085 ;
        RECT 15.780 87.360 18.455 87.915 ;
        RECT 24.740 87.520 26.840 88.120 ;
        RECT 16.115 87.205 18.455 87.360 ;
        RECT 24.140 87.220 25.340 87.520 ;
        RECT 26.240 87.220 27.140 87.520 ;
        RECT 16.115 86.635 18.810 87.205 ;
        RECT 24.140 86.920 25.640 87.220 ;
        RECT 25.940 86.920 27.740 87.220 ;
        RECT 16.455 86.495 18.810 86.635 ;
        RECT 23.840 86.620 24.440 86.920 ;
        RECT 25.040 86.620 26.540 86.920 ;
        RECT 27.140 86.620 27.740 86.920 ;
        RECT 16.455 85.915 19.170 86.495 ;
        RECT 23.840 86.320 24.140 86.620 ;
        RECT 16.810 85.790 19.170 85.915 ;
        RECT 23.540 86.020 24.140 86.320 ;
        RECT 16.810 85.205 19.540 85.790 ;
        RECT 17.170 85.090 19.540 85.205 ;
        RECT 23.540 85.720 24.440 86.020 ;
        RECT 25.340 85.720 26.240 86.620 ;
        RECT 27.440 86.320 27.740 86.620 ;
        RECT 38.110 86.420 38.560 89.465 ;
        RECT 39.465 89.180 42.345 89.465 ;
        RECT 39.465 88.925 42.800 89.180 ;
        RECT 39.900 88.615 42.800 88.925 ;
        RECT 50.910 88.740 59.750 90.950 ;
        RECT 88.480 88.740 97.320 90.950 ;
        RECT 107.840 91.470 111.055 91.520 ;
        RECT 107.840 90.925 119.630 91.470 ;
        RECT 107.415 90.910 119.630 90.925 ;
        RECT 107.415 90.740 110.660 90.910 ;
        RECT 107.415 90.335 110.255 90.740 ;
        RECT 106.980 90.125 110.255 90.335 ;
        RECT 106.980 89.755 109.840 90.125 ;
        RECT 106.535 89.520 109.840 89.755 ;
        RECT 106.535 89.180 109.415 89.520 ;
        RECT 39.900 88.335 43.270 88.615 ;
        RECT 40.345 88.060 43.270 88.335 ;
        RECT 40.345 87.755 43.745 88.060 ;
        RECT 40.800 87.510 43.745 87.755 ;
        RECT 40.800 87.180 44.230 87.510 ;
        RECT 41.270 86.970 44.230 87.180 ;
        RECT 41.270 86.615 44.725 86.970 ;
        RECT 27.440 86.020 28.040 86.320 ;
        RECT 27.140 85.720 28.040 86.020 ;
        RECT 17.170 84.495 19.920 85.090 ;
        RECT 23.540 84.520 28.040 85.720 ;
        RECT 29.550 85.860 38.560 86.420 ;
        RECT 41.745 86.435 44.725 86.615 ;
        RECT 50.910 86.530 57.540 88.740 ;
        RECT 90.690 86.530 97.320 88.740 ;
        RECT 106.080 88.925 109.415 89.180 ;
        RECT 114.750 89.250 117.150 89.550 ;
        RECT 114.750 88.950 117.450 89.250 ;
        RECT 106.080 88.615 108.980 88.925 ;
        RECT 105.610 88.335 108.980 88.615 ;
        RECT 114.150 88.350 118.050 88.950 ;
        RECT 119.070 88.550 119.630 90.910 ;
        RECT 123.290 91.370 123.890 91.670 ;
        RECT 123.290 91.070 124.190 91.370 ;
        RECT 125.090 91.070 125.990 91.970 ;
        RECT 127.190 91.670 127.490 91.970 ;
        RECT 132.350 91.775 134.915 92.290 ;
        RECT 127.190 91.370 127.790 91.670 ;
        RECT 132.350 91.550 134.635 91.775 ;
        RECT 126.890 91.070 127.790 91.370 ;
        RECT 123.290 89.870 127.790 91.070 ;
        RECT 132.050 91.030 134.635 91.550 ;
        RECT 132.050 90.815 134.350 91.030 ;
        RECT 131.745 90.290 134.350 90.815 ;
        RECT 131.745 90.085 134.050 90.290 ;
        RECT 123.590 89.270 127.490 89.870 ;
        RECT 124.190 88.970 126.890 89.270 ;
        RECT 124.190 88.670 126.590 88.970 ;
        RECT 128.620 88.750 129.070 89.740 ;
        RECT 131.425 89.550 134.050 90.085 ;
        RECT 131.425 89.360 133.745 89.550 ;
        RECT 131.100 88.815 133.745 89.360 ;
        RECT 131.100 88.750 133.425 88.815 ;
        RECT 105.610 88.060 108.535 88.335 ;
        RECT 105.135 87.755 108.535 88.060 ;
        RECT 105.135 87.510 108.080 87.755 ;
        RECT 104.650 87.180 108.080 87.510 ;
        RECT 104.650 86.970 107.610 87.180 ;
        RECT 104.155 86.615 107.610 86.970 ;
        RECT 113.850 87.150 118.350 88.350 ;
        RECT 128.620 88.300 133.425 88.750 ;
        RECT 130.765 88.085 133.425 88.300 ;
        RECT 130.765 87.915 133.100 88.085 ;
        RECT 130.425 87.360 133.100 87.915 ;
        RECT 130.425 87.205 132.765 87.360 ;
        RECT 130.110 87.190 132.765 87.205 ;
        RECT 113.850 86.850 114.750 87.150 ;
        RECT 41.745 86.060 45.230 86.435 ;
        RECT 17.540 84.395 19.920 84.495 ;
        RECT 17.540 83.790 20.310 84.395 ;
        RECT 23.840 83.920 27.740 84.520 ;
        RECT 17.920 83.705 20.310 83.790 ;
        RECT 17.920 83.090 20.705 83.705 ;
        RECT 24.440 83.620 27.140 83.920 ;
        RECT 28.760 83.820 29.320 84.320 ;
        RECT 29.550 83.820 30.110 85.860 ;
        RECT 38.110 85.370 38.560 85.860 ;
        RECT 42.230 85.915 45.230 86.060 ;
        RECT 42.230 85.510 45.745 85.915 ;
        RECT 33.680 84.680 36.080 84.980 ;
        RECT 33.680 84.380 36.380 84.680 ;
        RECT 24.440 83.320 26.840 83.620 ;
        RECT 18.310 83.020 20.705 83.090 ;
        RECT 28.760 83.260 30.110 83.820 ;
        RECT 33.080 83.780 36.980 84.380 ;
        RECT 38.000 83.980 38.560 85.370 ;
        RECT 42.725 85.400 45.745 85.510 ;
        RECT 42.725 84.970 46.265 85.400 ;
        RECT 43.230 84.895 46.265 84.970 ;
        RECT 43.230 84.435 46.800 84.895 ;
        RECT 43.745 84.400 46.800 84.435 ;
        RECT 43.745 83.915 47.340 84.400 ;
        RECT 53.120 84.320 55.330 86.530 ;
        RECT 92.900 84.320 95.110 86.530 ;
        RECT 104.155 86.435 107.135 86.615 ;
        RECT 113.850 86.550 114.450 86.850 ;
        RECT 103.650 86.060 107.135 86.435 ;
        RECT 114.150 86.250 114.450 86.550 ;
        RECT 115.650 86.250 116.550 87.150 ;
        RECT 117.450 86.850 118.350 87.150 ;
        RECT 117.750 86.550 118.350 86.850 ;
        RECT 130.070 86.635 132.765 87.190 ;
        RECT 117.750 86.250 118.050 86.550 ;
        RECT 130.070 86.495 132.425 86.635 ;
        RECT 103.650 85.915 106.650 86.060 ;
        RECT 114.150 85.950 114.750 86.250 ;
        RECT 115.350 85.950 116.850 86.250 ;
        RECT 117.450 85.950 118.050 86.250 ;
        RECT 103.135 85.510 106.650 85.915 ;
        RECT 114.450 85.650 115.950 85.950 ;
        RECT 116.250 85.650 118.050 85.950 ;
        RECT 129.710 85.915 132.425 86.495 ;
        RECT 129.710 85.790 132.070 85.915 ;
        RECT 103.135 85.400 106.155 85.510 ;
        RECT 102.615 84.970 106.155 85.400 ;
        RECT 114.450 85.350 115.650 85.650 ;
        RECT 116.550 85.350 117.450 85.650 ;
        RECT 102.615 84.895 105.650 84.970 ;
        RECT 102.080 84.495 105.650 84.895 ;
        RECT 115.050 84.750 117.150 85.350 ;
        RECT 129.340 85.205 132.070 85.790 ;
        RECT 129.340 85.090 131.710 85.205 ;
        RECT 102.080 84.400 109.090 84.495 ;
        RECT 113.250 84.450 113.550 84.750 ;
        RECT 115.050 84.450 115.350 84.750 ;
        RECT 115.650 84.450 115.950 84.750 ;
        RECT 116.250 84.450 116.550 84.750 ;
        RECT 116.850 84.450 117.150 84.750 ;
        RECT 118.650 84.450 118.950 84.750 ;
        RECT 128.960 84.495 131.710 85.090 ;
        RECT 101.540 84.045 109.090 84.400 ;
        RECT 101.540 83.915 105.135 84.045 ;
        RECT 18.310 82.395 21.110 83.020 ;
        RECT 28.760 82.930 29.320 83.260 ;
        RECT 18.705 82.335 21.110 82.395 ;
        RECT 32.780 82.580 37.280 83.780 ;
        RECT 44.265 83.440 47.890 83.915 ;
        RECT 100.990 83.440 104.615 83.915 ;
        RECT 44.265 83.400 48.445 83.440 ;
        RECT 44.800 82.970 48.445 83.400 ;
        RECT 100.435 83.400 104.615 83.440 ;
        RECT 100.435 82.970 104.080 83.400 ;
        RECT 44.800 82.895 49.010 82.970 ;
        RECT 18.705 81.705 21.525 82.335 ;
        RECT 32.780 82.280 33.680 82.580 ;
        RECT 32.780 81.980 33.380 82.280 ;
        RECT 19.110 81.665 21.525 81.705 ;
        RECT 33.080 81.680 33.380 81.980 ;
        RECT 34.580 81.680 35.480 82.580 ;
        RECT 36.380 82.280 37.280 82.580 ;
        RECT 45.340 82.515 49.010 82.895 ;
        RECT 99.870 82.895 104.080 82.970 ;
        RECT 99.870 82.515 103.540 82.895 ;
        RECT 45.340 82.400 49.585 82.515 ;
        RECT 36.680 81.980 37.280 82.280 ;
        RECT 45.890 82.070 49.585 82.400 ;
        RECT 99.295 82.400 103.540 82.515 ;
        RECT 99.295 82.070 102.990 82.400 ;
        RECT 36.680 81.680 36.980 81.980 ;
        RECT 45.890 81.915 50.165 82.070 ;
        RECT 19.110 81.020 21.945 81.665 ;
        RECT 33.080 81.380 33.680 81.680 ;
        RECT 34.280 81.380 35.780 81.680 ;
        RECT 36.380 81.380 36.980 81.680 ;
        RECT 46.445 81.635 50.165 81.915 ;
        RECT 98.715 81.915 102.990 82.070 ;
        RECT 98.715 81.635 102.435 81.915 ;
        RECT 46.445 81.440 50.755 81.635 ;
        RECT 19.525 80.995 21.945 81.020 ;
        RECT 33.380 81.080 34.880 81.380 ;
        RECT 35.180 81.080 36.980 81.380 ;
        RECT 47.010 81.210 50.755 81.440 ;
        RECT 98.125 81.440 102.435 81.635 ;
        RECT 98.125 81.210 101.870 81.440 ;
        RECT 19.525 80.335 22.375 80.995 ;
        RECT 33.380 80.780 34.580 81.080 ;
        RECT 35.480 80.780 36.380 81.080 ;
        RECT 47.010 80.970 51.350 81.210 ;
        RECT 47.585 80.795 51.350 80.970 ;
        RECT 97.530 80.970 101.870 81.210 ;
        RECT 97.530 80.795 101.295 80.970 ;
        RECT 19.945 80.330 22.375 80.335 ;
        RECT 19.945 79.670 22.815 80.330 ;
        RECT 33.980 80.180 36.080 80.780 ;
        RECT 47.585 80.515 51.955 80.795 ;
        RECT 48.165 80.390 51.955 80.515 ;
        RECT 96.925 80.515 101.295 80.795 ;
        RECT 96.925 80.390 100.715 80.515 ;
        RECT 32.180 79.880 32.480 80.180 ;
        RECT 33.980 79.880 34.280 80.180 ;
        RECT 34.580 79.880 34.880 80.180 ;
        RECT 35.180 79.880 35.480 80.180 ;
        RECT 35.780 79.880 36.080 80.180 ;
        RECT 37.580 79.880 37.880 80.180 ;
        RECT 48.165 80.070 52.570 80.390 ;
        RECT 48.755 79.995 52.570 80.070 ;
        RECT 96.310 80.070 100.715 80.390 ;
        RECT 108.640 80.080 109.090 84.045 ;
        RECT 112.950 84.150 113.850 84.450 ;
        RECT 118.350 84.150 119.250 84.450 ;
        RECT 128.960 84.395 131.340 84.495 ;
        RECT 112.950 83.850 114.150 84.150 ;
        RECT 118.050 83.850 119.250 84.150 ;
        RECT 112.950 83.550 114.750 83.850 ;
        RECT 117.450 83.550 119.250 83.850 ;
        RECT 128.570 83.790 131.340 84.395 ;
        RECT 128.570 83.705 130.960 83.790 ;
        RECT 112.950 83.250 115.350 83.550 ;
        RECT 116.850 83.250 118.950 83.550 ;
        RECT 114.750 82.950 115.950 83.250 ;
        RECT 116.250 82.950 117.450 83.250 ;
        RECT 128.175 83.090 130.960 83.705 ;
        RECT 128.175 83.020 130.570 83.090 ;
        RECT 115.350 82.350 116.850 82.950 ;
        RECT 127.770 82.395 130.570 83.020 ;
        RECT 114.750 82.050 115.950 82.350 ;
        RECT 116.250 82.050 117.450 82.350 ;
        RECT 127.770 82.335 130.175 82.395 ;
        RECT 114.150 81.750 115.350 82.050 ;
        RECT 116.850 81.750 118.050 82.050 ;
        RECT 113.250 81.450 115.050 81.750 ;
        RECT 117.150 81.450 118.950 81.750 ;
        RECT 127.355 81.705 130.175 82.335 ;
        RECT 127.355 81.665 129.770 81.705 ;
        RECT 112.950 80.850 114.450 81.450 ;
        RECT 117.750 80.850 119.250 81.450 ;
        RECT 126.935 81.020 129.770 81.665 ;
        RECT 126.935 80.995 129.355 81.020 ;
        RECT 113.250 80.550 114.150 80.850 ;
        RECT 115.050 80.550 115.350 80.850 ;
        RECT 115.650 80.550 115.950 80.850 ;
        RECT 116.250 80.550 116.550 80.850 ;
        RECT 116.850 80.550 117.150 80.850 ;
        RECT 118.050 80.550 118.950 80.850 ;
        RECT 96.310 79.995 100.125 80.070 ;
        RECT 19.945 79.665 23.265 79.670 ;
        RECT 20.375 79.015 23.265 79.665 ;
        RECT 31.880 79.580 32.780 79.880 ;
        RECT 37.280 79.580 38.180 79.880 ;
        RECT 48.755 79.635 53.185 79.995 ;
        RECT 31.880 79.280 33.080 79.580 ;
        RECT 36.980 79.280 38.180 79.580 ;
        RECT 20.375 78.995 23.720 79.015 ;
        RECT 20.815 78.370 23.720 78.995 ;
        RECT 31.880 78.980 33.680 79.280 ;
        RECT 36.380 78.980 38.180 79.280 ;
        RECT 49.350 79.610 53.185 79.635 ;
        RECT 95.695 79.635 100.125 79.995 ;
        RECT 95.695 79.610 99.530 79.635 ;
        RECT 49.350 79.240 53.810 79.610 ;
        RECT 95.070 79.240 99.530 79.610 ;
        RECT 49.350 79.210 54.440 79.240 ;
        RECT 31.880 78.680 34.280 78.980 ;
        RECT 35.780 78.680 37.880 78.980 ;
        RECT 49.955 78.880 54.440 79.210 ;
        RECT 94.440 79.210 99.530 79.240 ;
        RECT 104.210 79.390 106.610 79.690 ;
        RECT 94.440 78.880 98.925 79.210 ;
        RECT 104.210 79.090 106.910 79.390 ;
        RECT 49.955 78.795 55.080 78.880 ;
        RECT 33.680 78.380 34.880 78.680 ;
        RECT 35.180 78.380 36.380 78.680 ;
        RECT 50.220 78.530 55.080 78.795 ;
        RECT 93.800 78.795 98.925 78.880 ;
        RECT 93.800 78.530 98.310 78.795 ;
        RECT 50.220 78.390 55.725 78.530 ;
        RECT 20.815 78.330 24.185 78.370 ;
        RECT 21.265 77.730 24.185 78.330 ;
        RECT 34.280 77.780 35.780 78.380 ;
        RECT 21.265 77.670 24.655 77.730 ;
        RECT 21.720 77.095 24.655 77.670 ;
        RECT 33.680 77.480 34.880 77.780 ;
        RECT 35.180 77.480 36.380 77.780 ;
        RECT 33.080 77.180 34.280 77.480 ;
        RECT 35.780 77.180 36.980 77.480 ;
        RECT 21.720 77.015 25.135 77.095 ;
        RECT 22.185 76.465 25.135 77.015 ;
        RECT 32.180 76.880 33.980 77.180 ;
        RECT 36.080 76.880 37.880 77.180 ;
        RECT 22.185 76.370 25.625 76.465 ;
        RECT 22.655 75.840 25.625 76.370 ;
        RECT 31.880 76.280 33.380 76.880 ;
        RECT 36.680 76.280 38.180 76.880 ;
        RECT 32.180 75.980 33.080 76.280 ;
        RECT 33.980 75.980 34.280 76.280 ;
        RECT 34.580 75.980 34.880 76.280 ;
        RECT 35.180 75.980 35.480 76.280 ;
        RECT 35.780 75.980 36.080 76.280 ;
        RECT 36.980 75.980 37.880 76.280 ;
        RECT 22.655 75.730 26.120 75.840 ;
        RECT 23.135 75.225 26.120 75.730 ;
        RECT 33.980 75.380 36.080 75.980 ;
        RECT 50.220 75.700 50.670 78.390 ;
        RECT 51.185 78.190 55.725 78.390 ;
        RECT 93.155 78.390 98.310 78.530 ;
        RECT 103.610 78.490 107.510 79.090 ;
        RECT 108.530 78.690 109.090 80.080 ;
        RECT 115.050 79.950 117.150 80.550 ;
        RECT 126.505 80.335 129.355 80.995 ;
        RECT 126.505 80.330 128.935 80.335 ;
        RECT 114.450 79.650 115.650 79.950 ;
        RECT 116.550 79.650 117.450 79.950 ;
        RECT 126.065 79.670 128.935 80.330 ;
        RECT 125.615 79.665 128.935 79.670 ;
        RECT 114.450 79.350 115.950 79.650 ;
        RECT 116.250 79.350 118.050 79.650 ;
        RECT 114.150 79.050 114.750 79.350 ;
        RECT 115.350 79.050 116.850 79.350 ;
        RECT 117.450 79.050 118.050 79.350 ;
        RECT 114.150 78.750 114.450 79.050 ;
        RECT 93.155 78.190 97.695 78.390 ;
        RECT 51.185 77.995 56.375 78.190 ;
        RECT 51.810 77.865 56.375 77.995 ;
        RECT 92.505 77.995 97.695 78.190 ;
        RECT 92.505 77.865 97.070 77.995 ;
        RECT 51.810 77.610 57.030 77.865 ;
        RECT 52.440 77.550 57.030 77.610 ;
        RECT 91.850 77.610 97.070 77.865 ;
        RECT 91.850 77.550 96.440 77.610 ;
        RECT 52.440 77.245 57.695 77.550 ;
        RECT 91.185 77.245 96.440 77.550 ;
        RECT 52.440 77.240 58.360 77.245 ;
        RECT 53.080 76.950 58.360 77.240 ;
        RECT 90.520 77.240 96.440 77.245 ;
        RECT 103.310 77.290 107.810 78.490 ;
        RECT 90.520 76.950 95.800 77.240 ;
        RECT 53.080 76.880 59.030 76.950 ;
        RECT 53.725 76.670 59.030 76.880 ;
        RECT 89.850 76.880 95.800 76.950 ;
        RECT 103.310 76.990 104.210 77.290 ;
        RECT 89.850 76.670 95.375 76.880 ;
        RECT 103.310 76.690 103.910 76.990 ;
        RECT 53.725 76.530 59.710 76.670 ;
        RECT 54.375 76.400 59.710 76.530 ;
        RECT 89.170 76.530 95.375 76.670 ;
        RECT 89.170 76.400 94.505 76.530 ;
        RECT 54.375 76.190 60.390 76.400 ;
        RECT 55.030 76.145 60.390 76.190 ;
        RECT 88.490 76.190 94.505 76.400 ;
        RECT 88.490 76.145 93.850 76.190 ;
        RECT 55.030 75.900 61.080 76.145 ;
        RECT 87.800 75.900 93.850 76.145 ;
        RECT 55.030 75.865 61.770 75.900 ;
        RECT 23.135 75.095 26.625 75.225 ;
        RECT 23.625 74.615 26.625 75.095 ;
        RECT 33.380 75.080 34.580 75.380 ;
        RECT 35.480 75.080 36.380 75.380 ;
        RECT 33.380 74.780 34.880 75.080 ;
        RECT 35.180 74.780 36.980 75.080 ;
        RECT 23.625 74.465 27.135 74.615 ;
        RECT 24.120 74.010 27.135 74.465 ;
        RECT 33.080 74.480 33.680 74.780 ;
        RECT 34.280 74.480 35.780 74.780 ;
        RECT 36.380 74.480 36.980 74.780 ;
        RECT 45.790 75.010 48.190 75.310 ;
        RECT 45.790 74.710 48.490 75.010 ;
        RECT 33.080 74.180 33.380 74.480 ;
        RECT 24.120 73.840 27.655 74.010 ;
        RECT 24.625 73.415 27.655 73.840 ;
        RECT 32.780 73.880 33.380 74.180 ;
        RECT 32.780 73.580 33.680 73.880 ;
        RECT 34.580 73.580 35.480 74.480 ;
        RECT 36.680 74.180 36.980 74.480 ;
        RECT 36.680 73.880 37.280 74.180 ;
        RECT 45.190 74.110 49.090 74.710 ;
        RECT 50.110 74.310 50.670 75.700 ;
        RECT 55.695 75.670 61.770 75.865 ;
        RECT 87.110 75.865 93.850 75.900 ;
        RECT 94.925 76.165 95.375 76.530 ;
        RECT 103.610 76.390 103.910 76.690 ;
        RECT 105.110 76.390 106.010 77.290 ;
        RECT 106.910 76.990 107.810 77.290 ;
        RECT 107.210 76.690 107.810 76.990 ;
        RECT 113.850 78.450 114.450 78.750 ;
        RECT 113.850 78.150 114.750 78.450 ;
        RECT 115.650 78.150 116.550 79.050 ;
        RECT 117.750 78.750 118.050 79.050 ;
        RECT 125.615 79.015 128.505 79.665 ;
        RECT 125.160 78.995 128.505 79.015 ;
        RECT 117.750 78.450 118.350 78.750 ;
        RECT 117.450 78.150 118.350 78.450 ;
        RECT 125.160 78.370 128.065 78.995 ;
        RECT 113.850 76.950 118.350 78.150 ;
        RECT 124.695 78.330 128.065 78.370 ;
        RECT 124.695 77.730 127.615 78.330 ;
        RECT 124.225 77.670 127.615 77.730 ;
        RECT 124.225 77.095 127.160 77.670 ;
        RECT 123.745 77.015 127.160 77.095 ;
        RECT 107.210 76.390 107.510 76.690 ;
        RECT 87.110 75.670 93.185 75.865 ;
        RECT 94.925 75.715 95.660 76.165 ;
        RECT 103.610 76.090 104.210 76.390 ;
        RECT 104.810 76.090 106.310 76.390 ;
        RECT 106.910 76.090 107.510 76.390 ;
        RECT 114.150 76.350 118.050 76.950 ;
        RECT 55.695 75.550 62.465 75.670 ;
        RECT 56.360 75.450 62.465 75.550 ;
        RECT 86.415 75.550 93.185 75.670 ;
        RECT 86.415 75.450 92.520 75.550 ;
        RECT 56.360 75.245 63.165 75.450 ;
        RECT 57.030 75.240 63.165 75.245 ;
        RECT 85.715 75.245 92.520 75.450 ;
        RECT 85.715 75.240 91.850 75.245 ;
        RECT 57.030 75.045 63.865 75.240 ;
        RECT 85.015 75.045 91.850 75.240 ;
        RECT 57.030 74.950 64.570 75.045 ;
        RECT 57.710 74.860 64.570 74.950 ;
        RECT 84.310 74.950 91.850 75.045 ;
        RECT 84.310 74.860 91.170 74.950 ;
        RECT 57.710 74.690 65.280 74.860 ;
        RECT 83.600 74.690 91.170 74.860 ;
        RECT 57.710 74.670 65.995 74.690 ;
        RECT 58.390 74.530 65.995 74.670 ;
        RECT 82.885 74.670 91.170 74.690 ;
        RECT 82.885 74.530 90.490 74.670 ;
        RECT 58.390 74.400 66.710 74.530 ;
        RECT 59.080 74.385 66.710 74.400 ;
        RECT 82.170 74.400 90.490 74.530 ;
        RECT 82.170 74.385 89.800 74.400 ;
        RECT 59.080 74.250 67.430 74.385 ;
        RECT 81.450 74.250 89.800 74.385 ;
        RECT 59.080 74.145 68.150 74.250 ;
        RECT 59.770 74.130 68.150 74.145 ;
        RECT 80.730 74.145 89.800 74.250 ;
        RECT 80.730 74.130 89.110 74.145 ;
        RECT 36.380 73.580 37.280 73.880 ;
        RECT 24.625 73.225 28.180 73.415 ;
        RECT 25.135 72.825 28.180 73.225 ;
        RECT 25.135 72.615 28.715 72.825 ;
        RECT 25.655 72.240 28.715 72.615 ;
        RECT 32.780 72.380 37.280 73.580 ;
        RECT 44.890 72.910 49.390 74.110 ;
        RECT 59.770 74.020 68.870 74.130 ;
        RECT 80.010 74.020 89.110 74.130 ;
        RECT 59.770 73.925 69.595 74.020 ;
        RECT 79.285 73.925 89.110 74.020 ;
        RECT 59.770 73.900 70.325 73.925 ;
        RECT 60.465 73.845 70.325 73.900 ;
        RECT 78.555 73.900 89.110 73.925 ;
        RECT 78.555 73.845 88.415 73.900 ;
        RECT 60.465 73.770 71.050 73.845 ;
        RECT 77.830 73.770 88.415 73.845 ;
        RECT 60.465 73.715 71.780 73.770 ;
        RECT 77.100 73.715 88.415 73.770 ;
        RECT 60.465 73.670 72.515 73.715 ;
        RECT 76.365 73.670 88.415 73.715 ;
        RECT 61.165 73.640 73.245 73.670 ;
        RECT 75.635 73.640 87.715 73.670 ;
        RECT 61.165 73.620 73.975 73.640 ;
        RECT 74.905 73.620 87.715 73.640 ;
        RECT 61.165 73.450 87.715 73.620 ;
        RECT 61.865 73.240 87.015 73.450 ;
        RECT 62.570 73.045 86.310 73.240 ;
        RECT 44.890 72.610 45.790 72.910 ;
        RECT 25.655 72.010 29.255 72.240 ;
        RECT 26.180 71.665 29.255 72.010 ;
        RECT 33.080 71.780 36.980 72.380 ;
        RECT 44.890 72.310 45.490 72.610 ;
        RECT 26.180 71.415 29.805 71.665 ;
        RECT 26.715 71.095 29.805 71.415 ;
        RECT 33.680 71.480 36.380 71.780 ;
        RECT 33.680 71.180 36.080 71.480 ;
        RECT 26.715 70.825 30.360 71.095 ;
        RECT 27.255 70.530 30.360 70.825 ;
        RECT 27.255 70.240 30.925 70.530 ;
        RECT 27.805 69.975 30.925 70.240 ;
        RECT 27.805 69.665 31.495 69.975 ;
        RECT 28.360 69.425 31.495 69.665 ;
        RECT 28.360 69.095 32.070 69.425 ;
        RECT 28.925 68.885 32.070 69.095 ;
        RECT 28.925 68.530 32.655 68.885 ;
        RECT 29.495 68.350 32.655 68.530 ;
        RECT 29.495 67.975 33.245 68.350 ;
        RECT 30.070 67.825 33.245 67.975 ;
        RECT 30.070 67.425 33.840 67.825 ;
        RECT 30.655 67.305 33.840 67.425 ;
        RECT 30.655 66.885 34.445 67.305 ;
        RECT 31.245 66.795 34.445 66.885 ;
        RECT 31.245 66.350 35.055 66.795 ;
        RECT 31.840 66.290 35.055 66.350 ;
        RECT 31.840 65.825 35.670 66.290 ;
        RECT 32.445 65.795 35.670 65.825 ;
        RECT 32.445 65.305 36.295 65.795 ;
        RECT 33.055 64.825 36.925 65.305 ;
        RECT 33.055 64.795 37.560 64.825 ;
        RECT 33.670 64.355 37.560 64.795 ;
        RECT 38.110 64.355 38.560 72.250 ;
        RECT 45.190 72.010 45.490 72.310 ;
        RECT 46.690 72.010 47.590 72.910 ;
        RECT 48.490 72.610 49.390 72.910 ;
        RECT 63.280 72.860 85.600 73.045 ;
        RECT 63.995 72.690 84.885 72.860 ;
        RECT 48.790 72.310 49.390 72.610 ;
        RECT 64.650 72.530 84.170 72.690 ;
        RECT 48.790 72.010 49.090 72.310 ;
        RECT 45.190 71.710 45.790 72.010 ;
        RECT 46.390 71.710 47.890 72.010 ;
        RECT 48.490 71.710 49.090 72.010 ;
        RECT 45.490 71.410 46.990 71.710 ;
        RECT 47.290 71.410 49.090 71.710 ;
        RECT 45.490 71.110 46.690 71.410 ;
        RECT 47.590 71.110 48.490 71.410 ;
        RECT 46.090 70.510 48.190 71.110 ;
        RECT 44.290 70.210 44.590 70.510 ;
        RECT 46.090 70.210 46.390 70.510 ;
        RECT 46.690 70.210 46.990 70.510 ;
        RECT 47.290 70.210 47.590 70.510 ;
        RECT 47.890 70.210 48.190 70.510 ;
        RECT 49.690 70.210 49.990 70.510 ;
        RECT 43.990 69.910 44.890 70.210 ;
        RECT 49.390 69.910 50.290 70.210 ;
        RECT 64.650 70.040 65.100 72.530 ;
        RECT 65.430 72.385 83.450 72.530 ;
        RECT 66.150 72.250 82.730 72.385 ;
        RECT 95.210 72.330 95.660 75.715 ;
        RECT 103.910 75.790 105.410 76.090 ;
        RECT 105.710 75.790 107.510 76.090 ;
        RECT 114.750 76.050 117.450 76.350 ;
        RECT 103.910 75.490 105.110 75.790 ;
        RECT 106.010 75.490 106.910 75.790 ;
        RECT 114.750 75.750 117.150 76.050 ;
        RECT 119.180 75.830 119.630 76.820 ;
        RECT 123.745 76.465 126.695 77.015 ;
        RECT 123.255 76.370 126.695 76.465 ;
        RECT 123.255 75.840 126.225 76.370 ;
        RECT 122.760 75.830 126.225 75.840 ;
        RECT 119.180 75.730 126.225 75.830 ;
        RECT 104.510 74.890 106.610 75.490 ;
        RECT 119.180 75.380 125.745 75.730 ;
        RECT 122.760 75.225 125.745 75.380 ;
        RECT 122.255 75.095 125.745 75.225 ;
        RECT 102.710 74.590 103.010 74.890 ;
        RECT 104.510 74.590 104.810 74.890 ;
        RECT 105.110 74.590 105.410 74.890 ;
        RECT 105.710 74.590 106.010 74.890 ;
        RECT 106.310 74.590 106.610 74.890 ;
        RECT 108.110 74.590 108.410 74.890 ;
        RECT 122.255 74.615 125.255 75.095 ;
        RECT 102.410 74.290 103.310 74.590 ;
        RECT 107.810 74.290 108.710 74.590 ;
        RECT 102.410 73.990 103.610 74.290 ;
        RECT 107.510 73.990 108.710 74.290 ;
        RECT 121.745 74.465 125.255 74.615 ;
        RECT 121.745 74.010 124.760 74.465 ;
        RECT 102.410 73.690 104.210 73.990 ;
        RECT 106.910 73.690 108.710 73.990 ;
        RECT 121.225 73.840 124.760 74.010 ;
        RECT 102.410 73.390 104.810 73.690 ;
        RECT 106.310 73.390 108.410 73.690 ;
        RECT 121.225 73.415 124.255 73.840 ;
        RECT 104.210 73.090 105.410 73.390 ;
        RECT 105.710 73.090 106.910 73.390 ;
        RECT 120.700 73.225 124.255 73.415 ;
        RECT 104.810 72.490 106.310 73.090 ;
        RECT 120.700 72.825 123.745 73.225 ;
        RECT 120.165 72.615 123.745 72.825 ;
        RECT 66.870 72.130 82.010 72.250 ;
        RECT 67.595 72.020 81.285 72.130 ;
        RECT 68.325 71.925 80.555 72.020 ;
        RECT 69.050 71.845 79.830 71.925 ;
        RECT 69.780 71.770 79.100 71.845 ;
        RECT 70.515 71.715 78.365 71.770 ;
        RECT 71.245 71.670 77.635 71.715 ;
        RECT 71.975 71.640 76.905 71.670 ;
        RECT 72.710 71.620 76.170 71.640 ;
        RECT 73.440 71.610 75.435 71.620 ;
        RECT 43.990 69.610 45.190 69.910 ;
        RECT 49.090 69.610 50.290 69.910 ;
        RECT 43.990 69.310 45.790 69.610 ;
        RECT 48.490 69.310 50.290 69.610 ;
        RECT 60.220 69.350 62.620 69.650 ;
        RECT 43.990 69.010 46.390 69.310 ;
        RECT 47.890 69.010 49.990 69.310 ;
        RECT 60.220 69.050 62.920 69.350 ;
        RECT 45.790 68.710 46.990 69.010 ;
        RECT 47.290 68.710 48.490 69.010 ;
        RECT 46.390 68.110 47.890 68.710 ;
        RECT 59.620 68.450 63.520 69.050 ;
        RECT 64.540 68.650 65.100 70.040 ;
        RECT 80.100 68.880 80.550 71.925 ;
        RECT 90.780 71.640 93.180 71.940 ;
        RECT 90.780 71.340 93.480 71.640 ;
        RECT 90.180 70.740 94.080 71.340 ;
        RECT 95.100 70.940 95.660 72.330 ;
        RECT 104.210 72.190 105.410 72.490 ;
        RECT 105.710 72.190 106.910 72.490 ;
        RECT 120.165 72.240 123.225 72.615 ;
        RECT 103.610 71.890 104.810 72.190 ;
        RECT 106.310 71.890 107.510 72.190 ;
        RECT 119.625 72.010 123.225 72.240 ;
        RECT 102.710 71.590 104.510 71.890 ;
        RECT 106.610 71.590 108.410 71.890 ;
        RECT 119.625 71.665 122.700 72.010 ;
        RECT 102.410 70.990 103.910 71.590 ;
        RECT 107.210 70.990 108.710 71.590 ;
        RECT 119.075 71.415 122.700 71.665 ;
        RECT 119.075 71.095 122.165 71.415 ;
        RECT 89.880 69.540 94.380 70.740 ;
        RECT 102.710 70.690 103.610 70.990 ;
        RECT 104.510 70.690 104.810 70.990 ;
        RECT 105.110 70.690 105.410 70.990 ;
        RECT 105.710 70.690 106.010 70.990 ;
        RECT 106.310 70.690 106.610 70.990 ;
        RECT 107.510 70.690 108.410 70.990 ;
        RECT 118.520 70.825 122.165 71.095 ;
        RECT 104.510 70.090 106.610 70.690 ;
        RECT 118.520 70.530 121.625 70.825 ;
        RECT 117.955 70.240 121.625 70.530 ;
        RECT 89.880 69.240 90.780 69.540 ;
        RECT 89.880 68.940 90.480 69.240 ;
        RECT 45.790 67.810 46.990 68.110 ;
        RECT 47.290 67.810 48.490 68.110 ;
        RECT 45.190 67.510 46.390 67.810 ;
        RECT 47.890 67.510 49.090 67.810 ;
        RECT 44.290 67.210 46.090 67.510 ;
        RECT 48.190 67.210 49.990 67.510 ;
        RECT 59.320 67.250 63.820 68.450 ;
        RECT 75.670 68.190 78.070 68.490 ;
        RECT 75.670 67.890 78.370 68.190 ;
        RECT 75.070 67.290 78.970 67.890 ;
        RECT 79.990 67.490 80.550 68.880 ;
        RECT 90.180 68.640 90.480 68.940 ;
        RECT 91.680 68.640 92.580 69.540 ;
        RECT 93.480 69.240 94.380 69.540 ;
        RECT 103.910 69.790 105.110 70.090 ;
        RECT 106.010 69.790 106.910 70.090 ;
        RECT 117.955 69.975 121.075 70.240 ;
        RECT 103.910 69.490 105.410 69.790 ;
        RECT 105.710 69.490 107.510 69.790 ;
        RECT 93.780 68.940 94.380 69.240 ;
        RECT 103.610 69.190 104.210 69.490 ;
        RECT 104.810 69.190 106.310 69.490 ;
        RECT 106.910 69.190 107.510 69.490 ;
        RECT 117.385 69.665 121.075 69.975 ;
        RECT 117.385 69.425 120.520 69.665 ;
        RECT 93.780 68.640 94.080 68.940 ;
        RECT 103.610 68.890 103.910 69.190 ;
        RECT 90.180 68.340 90.780 68.640 ;
        RECT 91.380 68.340 92.880 68.640 ;
        RECT 93.480 68.340 94.080 68.640 ;
        RECT 90.480 68.040 91.980 68.340 ;
        RECT 92.280 68.040 94.080 68.340 ;
        RECT 103.310 68.590 103.910 68.890 ;
        RECT 103.310 68.290 104.210 68.590 ;
        RECT 105.110 68.290 106.010 69.190 ;
        RECT 107.210 68.890 107.510 69.190 ;
        RECT 116.810 69.095 120.520 69.425 ;
        RECT 107.210 68.590 107.810 68.890 ;
        RECT 116.810 68.885 119.955 69.095 ;
        RECT 106.910 68.290 107.810 68.590 ;
        RECT 116.225 68.530 119.955 68.885 ;
        RECT 116.225 68.350 119.385 68.530 ;
        RECT 90.480 67.740 91.680 68.040 ;
        RECT 92.580 67.740 93.480 68.040 ;
        RECT 43.990 66.610 45.490 67.210 ;
        RECT 48.790 66.610 50.290 67.210 ;
        RECT 59.320 66.950 60.220 67.250 ;
        RECT 59.320 66.650 59.920 66.950 ;
        RECT 44.290 66.310 45.190 66.610 ;
        RECT 46.090 66.310 46.390 66.610 ;
        RECT 46.690 66.310 46.990 66.610 ;
        RECT 47.290 66.310 47.590 66.610 ;
        RECT 47.890 66.310 48.190 66.610 ;
        RECT 49.090 66.310 49.990 66.610 ;
        RECT 59.620 66.350 59.920 66.650 ;
        RECT 61.120 66.350 62.020 67.250 ;
        RECT 62.920 66.950 63.820 67.250 ;
        RECT 63.220 66.650 63.820 66.950 ;
        RECT 63.220 66.350 63.520 66.650 ;
        RECT 46.090 65.710 48.190 66.310 ;
        RECT 59.620 66.050 60.220 66.350 ;
        RECT 60.820 66.050 62.320 66.350 ;
        RECT 62.920 66.050 63.520 66.350 ;
        RECT 59.920 65.750 61.420 66.050 ;
        RECT 61.720 65.750 63.520 66.050 ;
        RECT 74.770 66.090 79.270 67.290 ;
        RECT 91.080 67.140 93.180 67.740 ;
        RECT 89.280 66.840 89.580 67.140 ;
        RECT 91.080 66.840 91.380 67.140 ;
        RECT 91.680 66.840 91.980 67.140 ;
        RECT 92.280 66.840 92.580 67.140 ;
        RECT 92.880 66.840 93.180 67.140 ;
        RECT 94.680 66.840 94.980 67.140 ;
        RECT 103.310 67.090 107.810 68.290 ;
        RECT 115.635 67.975 119.385 68.350 ;
        RECT 115.635 67.825 118.810 67.975 ;
        RECT 115.040 67.425 118.810 67.825 ;
        RECT 115.040 67.305 118.225 67.425 ;
        RECT 74.770 65.790 75.670 66.090 ;
        RECT 45.490 65.410 46.690 65.710 ;
        RECT 47.590 65.410 48.490 65.710 ;
        RECT 59.920 65.450 61.120 65.750 ;
        RECT 62.020 65.450 62.920 65.750 ;
        RECT 74.770 65.490 75.370 65.790 ;
        RECT 45.490 65.110 46.990 65.410 ;
        RECT 47.290 65.110 49.090 65.410 ;
        RECT 45.190 64.810 45.790 65.110 ;
        RECT 46.390 64.810 47.890 65.110 ;
        RECT 48.490 64.810 49.090 65.110 ;
        RECT 60.520 64.850 62.620 65.450 ;
        RECT 75.070 65.190 75.370 65.490 ;
        RECT 76.570 65.190 77.470 66.090 ;
        RECT 78.370 65.790 79.270 66.090 ;
        RECT 78.670 65.490 79.270 65.790 ;
        RECT 88.980 66.540 89.880 66.840 ;
        RECT 94.380 66.540 95.280 66.840 ;
        RECT 88.980 66.240 90.180 66.540 ;
        RECT 94.080 66.240 95.280 66.540 ;
        RECT 103.610 66.490 107.510 67.090 ;
        RECT 88.980 65.940 90.780 66.240 ;
        RECT 93.480 65.940 95.280 66.240 ;
        RECT 104.210 66.190 106.910 66.490 ;
        RECT 88.980 65.640 91.380 65.940 ;
        RECT 92.880 65.640 94.980 65.940 ;
        RECT 104.210 65.890 106.610 66.190 ;
        RECT 78.670 65.190 78.970 65.490 ;
        RECT 90.780 65.340 91.980 65.640 ;
        RECT 92.280 65.340 93.480 65.640 ;
        RECT 75.070 64.890 75.670 65.190 ;
        RECT 76.270 64.890 77.770 65.190 ;
        RECT 78.370 64.890 78.970 65.190 ;
        RECT 45.190 64.510 45.490 64.810 ;
        RECT 33.670 64.290 38.560 64.355 ;
        RECT 34.295 63.890 38.560 64.290 ;
        RECT 44.890 64.210 45.490 64.510 ;
        RECT 44.890 63.910 45.790 64.210 ;
        RECT 46.690 63.910 47.590 64.810 ;
        RECT 48.790 64.510 49.090 64.810 ;
        RECT 58.720 64.550 59.020 64.850 ;
        RECT 60.520 64.550 60.820 64.850 ;
        RECT 61.120 64.550 61.420 64.850 ;
        RECT 61.720 64.550 62.020 64.850 ;
        RECT 62.320 64.550 62.620 64.850 ;
        RECT 64.120 64.550 64.420 64.850 ;
        RECT 75.370 64.590 76.870 64.890 ;
        RECT 77.170 64.590 78.970 64.890 ;
        RECT 91.380 64.740 92.880 65.340 ;
        RECT 48.790 64.210 49.390 64.510 ;
        RECT 48.490 63.910 49.390 64.210 ;
        RECT 34.295 63.795 38.845 63.890 ;
        RECT 34.925 63.435 38.845 63.795 ;
        RECT 34.925 63.305 39.500 63.435 ;
        RECT 35.560 62.985 39.500 63.305 ;
        RECT 35.560 62.825 40.160 62.985 ;
        RECT 36.200 62.545 40.160 62.825 ;
        RECT 44.890 62.710 49.390 63.910 ;
        RECT 58.420 64.250 59.320 64.550 ;
        RECT 63.820 64.250 64.720 64.550 ;
        RECT 75.370 64.290 76.570 64.590 ;
        RECT 77.470 64.290 78.370 64.590 ;
        RECT 90.780 64.440 91.980 64.740 ;
        RECT 92.280 64.440 93.480 64.740 ;
        RECT 58.420 63.950 59.620 64.250 ;
        RECT 63.520 63.950 64.720 64.250 ;
        RECT 58.420 63.650 60.220 63.950 ;
        RECT 62.920 63.650 64.720 63.950 ;
        RECT 75.970 63.690 78.070 64.290 ;
        RECT 90.180 64.140 91.380 64.440 ;
        RECT 92.880 64.140 94.080 64.440 ;
        RECT 89.280 63.840 91.080 64.140 ;
        RECT 93.180 63.840 94.980 64.140 ;
        RECT 58.420 63.350 60.820 63.650 ;
        RECT 62.320 63.350 64.420 63.650 ;
        RECT 74.170 63.390 74.470 63.690 ;
        RECT 75.970 63.390 76.270 63.690 ;
        RECT 76.570 63.390 76.870 63.690 ;
        RECT 77.170 63.390 77.470 63.690 ;
        RECT 77.770 63.390 78.070 63.690 ;
        RECT 79.570 63.390 79.870 63.690 ;
        RECT 60.220 63.050 61.420 63.350 ;
        RECT 61.720 63.050 62.920 63.350 ;
        RECT 73.870 63.090 74.770 63.390 ;
        RECT 79.270 63.090 80.170 63.390 ;
        RECT 88.980 63.240 90.480 63.840 ;
        RECT 93.780 63.240 95.280 63.840 ;
        RECT 36.200 62.355 40.825 62.545 ;
        RECT 36.845 62.115 40.825 62.355 ;
        RECT 36.845 61.890 41.495 62.115 ;
        RECT 45.190 62.110 49.090 62.710 ;
        RECT 37.500 61.695 41.495 61.890 ;
        RECT 45.790 61.810 48.490 62.110 ;
        RECT 37.500 61.435 42.165 61.695 ;
        RECT 45.790 61.510 48.190 61.810 ;
        RECT 38.160 61.280 42.165 61.435 ;
        RECT 38.160 60.985 42.850 61.280 ;
        RECT 38.825 60.875 42.850 60.985 ;
        RECT 38.825 60.545 43.535 60.875 ;
        RECT 39.495 60.480 43.535 60.545 ;
        RECT 39.495 60.115 44.225 60.480 ;
        RECT 40.165 60.090 44.225 60.115 ;
        RECT 40.165 59.710 44.920 60.090 ;
        RECT 40.165 59.695 45.620 59.710 ;
        RECT 40.850 59.340 45.620 59.695 ;
        RECT 40.850 59.280 46.325 59.340 ;
        RECT 41.535 58.980 46.325 59.280 ;
        RECT 41.535 58.875 47.035 58.980 ;
        RECT 42.225 58.625 47.035 58.875 ;
        RECT 42.225 58.480 47.745 58.625 ;
        RECT 42.920 58.285 47.745 58.480 ;
        RECT 42.920 58.090 48.465 58.285 ;
        RECT 43.620 57.950 48.465 58.090 ;
        RECT 43.620 57.710 49.190 57.950 ;
        RECT 44.325 57.625 49.190 57.710 ;
        RECT 44.325 57.340 49.915 57.625 ;
        RECT 45.035 57.305 49.915 57.340 ;
        RECT 50.220 57.305 50.670 62.580 ;
        RECT 60.820 62.450 62.320 63.050 ;
        RECT 73.870 62.790 75.070 63.090 ;
        RECT 78.970 62.790 80.170 63.090 ;
        RECT 89.280 62.940 90.180 63.240 ;
        RECT 91.080 62.940 91.380 63.240 ;
        RECT 91.680 62.940 91.980 63.240 ;
        RECT 92.280 62.940 92.580 63.240 ;
        RECT 92.880 62.940 93.180 63.240 ;
        RECT 94.080 62.940 94.980 63.240 ;
        RECT 108.640 62.985 109.090 66.960 ;
        RECT 114.435 66.885 118.225 67.305 ;
        RECT 114.435 66.795 117.635 66.885 ;
        RECT 113.825 66.350 117.635 66.795 ;
        RECT 113.825 66.290 117.040 66.350 ;
        RECT 113.210 65.825 117.040 66.290 ;
        RECT 113.210 65.795 116.435 65.825 ;
        RECT 112.585 65.305 116.435 65.795 ;
        RECT 111.955 64.825 115.825 65.305 ;
        RECT 111.320 64.795 115.825 64.825 ;
        RECT 111.320 64.355 115.210 64.795 ;
        RECT 110.680 64.290 115.210 64.355 ;
        RECT 110.680 63.890 114.585 64.290 ;
        RECT 110.035 63.795 114.585 63.890 ;
        RECT 110.035 63.435 113.955 63.795 ;
        RECT 109.380 63.305 113.955 63.435 ;
        RECT 109.380 62.985 113.320 63.305 ;
        RECT 73.870 62.490 75.670 62.790 ;
        RECT 78.370 62.490 80.170 62.790 ;
        RECT 60.220 62.150 61.420 62.450 ;
        RECT 61.720 62.150 62.920 62.450 ;
        RECT 73.870 62.190 76.270 62.490 ;
        RECT 77.770 62.190 79.870 62.490 ;
        RECT 91.080 62.340 93.180 62.940 ;
        RECT 108.640 62.825 113.320 62.985 ;
        RECT 108.640 62.545 112.680 62.825 ;
        RECT 108.055 62.355 112.680 62.545 ;
        RECT 59.620 61.850 60.820 62.150 ;
        RECT 62.320 61.850 63.520 62.150 ;
        RECT 75.670 61.890 76.870 62.190 ;
        RECT 77.170 61.890 78.370 62.190 ;
        RECT 90.480 62.040 91.680 62.340 ;
        RECT 92.580 62.040 93.480 62.340 ;
        RECT 108.055 62.115 112.035 62.355 ;
        RECT 58.720 61.550 60.520 61.850 ;
        RECT 62.620 61.550 64.420 61.850 ;
        RECT 58.420 60.950 59.920 61.550 ;
        RECT 63.220 60.950 64.720 61.550 ;
        RECT 76.270 61.290 77.770 61.890 ;
        RECT 90.480 61.740 91.980 62.040 ;
        RECT 92.280 61.740 94.080 62.040 ;
        RECT 90.180 61.440 90.780 61.740 ;
        RECT 91.380 61.440 92.880 61.740 ;
        RECT 93.480 61.440 94.080 61.740 ;
        RECT 107.385 61.890 112.035 62.115 ;
        RECT 107.385 61.695 111.380 61.890 ;
        RECT 75.670 60.990 76.870 61.290 ;
        RECT 77.170 60.990 78.370 61.290 ;
        RECT 90.180 61.140 90.480 61.440 ;
        RECT 58.720 60.650 59.620 60.950 ;
        RECT 60.520 60.650 60.820 60.950 ;
        RECT 61.120 60.650 61.420 60.950 ;
        RECT 61.720 60.650 62.020 60.950 ;
        RECT 62.320 60.650 62.620 60.950 ;
        RECT 63.520 60.650 64.420 60.950 ;
        RECT 75.070 60.690 76.270 60.990 ;
        RECT 77.770 60.690 78.970 60.990 ;
        RECT 89.880 60.840 90.480 61.140 ;
        RECT 60.520 60.050 62.620 60.650 ;
        RECT 74.170 60.390 75.970 60.690 ;
        RECT 78.070 60.390 79.870 60.690 ;
        RECT 89.880 60.540 90.780 60.840 ;
        RECT 91.680 60.540 92.580 61.440 ;
        RECT 93.780 61.140 94.080 61.440 ;
        RECT 106.715 61.435 111.380 61.695 ;
        RECT 106.715 61.280 110.720 61.435 ;
        RECT 93.780 60.840 94.380 61.140 ;
        RECT 106.030 60.985 110.720 61.280 ;
        RECT 106.030 60.875 110.055 60.985 ;
        RECT 93.480 60.540 94.380 60.840 ;
        RECT 59.920 59.750 61.120 60.050 ;
        RECT 62.020 59.750 62.920 60.050 ;
        RECT 73.870 59.790 75.370 60.390 ;
        RECT 78.670 59.790 80.170 60.390 ;
        RECT 59.920 59.450 61.420 59.750 ;
        RECT 61.720 59.450 63.520 59.750 ;
        RECT 74.170 59.490 75.070 59.790 ;
        RECT 75.970 59.490 76.270 59.790 ;
        RECT 76.570 59.490 76.870 59.790 ;
        RECT 77.170 59.490 77.470 59.790 ;
        RECT 77.770 59.490 78.070 59.790 ;
        RECT 78.970 59.490 79.870 59.790 ;
        RECT 59.620 59.150 60.220 59.450 ;
        RECT 60.820 59.150 62.320 59.450 ;
        RECT 62.920 59.150 63.520 59.450 ;
        RECT 59.620 58.850 59.920 59.150 ;
        RECT 45.035 57.000 50.670 57.305 ;
        RECT 59.320 58.550 59.920 58.850 ;
        RECT 59.320 58.250 60.220 58.550 ;
        RECT 61.120 58.250 62.020 59.150 ;
        RECT 63.220 58.850 63.520 59.150 ;
        RECT 75.970 58.890 78.070 59.490 ;
        RECT 89.880 59.340 94.380 60.540 ;
        RECT 105.345 60.545 110.055 60.875 ;
        RECT 105.345 60.480 109.385 60.545 ;
        RECT 104.655 60.115 109.385 60.480 ;
        RECT 104.655 60.090 108.715 60.115 ;
        RECT 103.960 59.710 108.715 60.090 ;
        RECT 103.260 59.695 108.715 59.710 ;
        RECT 103.260 59.340 108.030 59.695 ;
        RECT 63.220 58.550 63.820 58.850 ;
        RECT 62.920 58.250 63.820 58.550 ;
        RECT 75.370 58.590 76.570 58.890 ;
        RECT 77.470 58.590 78.370 58.890 ;
        RECT 90.180 58.740 94.080 59.340 ;
        RECT 102.555 59.280 108.030 59.340 ;
        RECT 75.370 58.290 76.870 58.590 ;
        RECT 77.170 58.290 78.970 58.590 ;
        RECT 59.320 57.050 63.820 58.250 ;
        RECT 75.070 57.990 75.670 58.290 ;
        RECT 76.270 57.990 77.770 58.290 ;
        RECT 78.370 57.990 78.970 58.290 ;
        RECT 90.780 58.440 93.480 58.740 ;
        RECT 90.780 58.140 93.180 58.440 ;
        RECT 75.070 57.690 75.370 57.990 ;
        RECT 74.770 57.390 75.370 57.690 ;
        RECT 74.770 57.090 75.670 57.390 ;
        RECT 76.570 57.090 77.470 57.990 ;
        RECT 78.670 57.690 78.970 57.990 ;
        RECT 78.670 57.390 79.270 57.690 ;
        RECT 78.370 57.090 79.270 57.390 ;
        RECT 45.035 56.980 51.380 57.000 ;
        RECT 45.745 56.700 51.380 56.980 ;
        RECT 45.745 56.625 52.120 56.700 ;
        RECT 46.465 56.415 52.120 56.625 ;
        RECT 59.620 56.450 63.520 57.050 ;
        RECT 46.465 56.285 52.860 56.415 ;
        RECT 47.190 56.135 52.860 56.285 ;
        RECT 60.220 56.150 62.920 56.450 ;
        RECT 47.190 55.950 53.605 56.135 ;
        RECT 47.915 55.865 53.605 55.950 ;
        RECT 47.915 55.625 54.355 55.865 ;
        RECT 60.220 55.850 62.620 56.150 ;
        RECT 48.645 55.605 54.355 55.625 ;
        RECT 48.645 55.355 55.110 55.605 ;
        RECT 48.645 55.305 55.865 55.355 ;
        RECT 49.380 55.110 55.865 55.305 ;
        RECT 49.380 55.000 56.620 55.110 ;
        RECT 50.120 54.880 56.620 55.000 ;
        RECT 50.120 54.700 57.385 54.880 ;
        RECT 50.860 54.660 57.385 54.700 ;
        RECT 50.860 54.445 58.150 54.660 ;
        RECT 50.860 54.415 58.915 54.445 ;
        RECT 51.605 54.245 58.915 54.415 ;
        RECT 51.605 54.135 59.685 54.245 ;
        RECT 52.355 54.050 59.685 54.135 ;
        RECT 52.355 53.865 60.460 54.050 ;
        RECT 53.110 53.695 61.235 53.865 ;
        RECT 53.110 53.605 62.010 53.695 ;
        RECT 53.865 53.530 62.010 53.605 ;
        RECT 53.865 53.375 62.790 53.530 ;
        RECT 53.865 53.355 63.570 53.375 ;
        RECT 54.620 53.230 63.570 53.355 ;
        RECT 54.620 53.110 64.355 53.230 ;
        RECT 55.385 53.095 64.355 53.110 ;
        RECT 64.650 53.095 65.100 56.920 ;
        RECT 74.770 55.890 79.270 57.090 ;
        RECT 95.210 56.135 95.660 59.210 ;
        RECT 102.555 58.980 107.345 59.280 ;
        RECT 101.845 58.875 107.345 58.980 ;
        RECT 101.845 58.625 106.655 58.875 ;
        RECT 101.135 58.480 106.655 58.625 ;
        RECT 101.135 58.285 105.960 58.480 ;
        RECT 100.415 58.090 105.960 58.285 ;
        RECT 100.415 57.950 105.260 58.090 ;
        RECT 99.690 57.710 105.260 57.950 ;
        RECT 99.690 57.625 104.555 57.710 ;
        RECT 98.965 57.340 104.555 57.625 ;
        RECT 98.965 57.305 103.845 57.340 ;
        RECT 98.235 57.000 103.845 57.305 ;
        RECT 97.500 56.980 103.845 57.000 ;
        RECT 97.500 56.700 103.135 56.980 ;
        RECT 96.760 56.625 103.135 56.700 ;
        RECT 96.760 56.415 102.415 56.625 ;
        RECT 96.020 56.285 102.415 56.415 ;
        RECT 96.020 56.135 101.690 56.285 ;
        RECT 95.210 55.950 101.690 56.135 ;
        RECT 75.070 55.290 78.970 55.890 ;
        RECT 95.210 55.865 100.965 55.950 ;
        RECT 75.670 54.990 78.370 55.290 ;
        RECT 75.670 54.690 78.070 54.990 ;
        RECT 55.385 52.970 65.140 53.095 ;
        RECT 80.100 53.065 80.550 55.760 ;
        RECT 94.525 55.625 100.965 55.865 ;
        RECT 94.525 55.605 100.235 55.625 ;
        RECT 93.770 55.355 100.235 55.605 ;
        RECT 93.015 55.305 100.235 55.355 ;
        RECT 93.015 55.110 99.500 55.305 ;
        RECT 92.260 55.000 99.500 55.110 ;
        RECT 92.260 54.880 98.760 55.000 ;
        RECT 91.495 54.700 98.760 54.880 ;
        RECT 91.495 54.660 98.020 54.700 ;
        RECT 90.730 54.445 98.020 54.660 ;
        RECT 89.965 54.415 98.020 54.445 ;
        RECT 89.965 54.245 97.275 54.415 ;
        RECT 89.195 54.135 97.275 54.245 ;
        RECT 89.195 54.050 96.525 54.135 ;
        RECT 88.420 53.865 96.525 54.050 ;
        RECT 87.645 53.695 95.770 53.865 ;
        RECT 86.870 53.605 95.770 53.695 ;
        RECT 86.870 53.530 95.015 53.605 ;
        RECT 86.090 53.375 95.015 53.530 ;
        RECT 85.310 53.355 95.015 53.375 ;
        RECT 85.310 53.230 94.260 53.355 ;
        RECT 84.525 53.110 94.260 53.230 ;
        RECT 84.525 53.095 93.495 53.110 ;
        RECT 55.385 52.880 65.925 52.970 ;
        RECT 56.150 52.855 65.925 52.880 ;
        RECT 56.150 52.750 66.710 52.855 ;
        RECT 56.150 52.660 67.500 52.750 ;
        RECT 56.915 52.655 67.500 52.660 ;
        RECT 80.100 52.655 80.825 53.065 ;
        RECT 83.740 52.970 93.495 53.095 ;
        RECT 82.955 52.880 93.495 52.970 ;
        RECT 82.955 52.855 92.730 52.880 ;
        RECT 82.170 52.750 92.730 52.855 ;
        RECT 81.380 52.660 92.730 52.750 ;
        RECT 81.380 52.655 91.965 52.660 ;
        RECT 56.915 52.570 68.290 52.655 ;
        RECT 80.100 52.570 91.965 52.655 ;
        RECT 56.915 52.495 69.085 52.570 ;
        RECT 79.795 52.495 91.965 52.570 ;
        RECT 56.915 52.445 69.875 52.495 ;
        RECT 57.685 52.435 69.875 52.445 ;
        RECT 79.005 52.445 91.965 52.495 ;
        RECT 79.005 52.435 91.195 52.445 ;
        RECT 57.685 52.380 70.670 52.435 ;
        RECT 78.210 52.380 91.195 52.435 ;
        RECT 57.685 52.335 71.465 52.380 ;
        RECT 77.415 52.335 91.195 52.380 ;
        RECT 57.685 52.300 72.260 52.335 ;
        RECT 76.620 52.300 91.195 52.335 ;
        RECT 57.685 52.275 73.055 52.300 ;
        RECT 75.825 52.275 91.195 52.300 ;
        RECT 57.685 52.260 73.850 52.275 ;
        RECT 75.030 52.260 91.195 52.275 ;
        RECT 57.685 52.245 91.195 52.260 ;
        RECT 58.460 52.050 90.420 52.245 ;
        RECT 59.235 51.865 89.645 52.050 ;
        RECT 60.010 51.695 88.870 51.865 ;
        RECT 60.790 51.530 88.090 51.695 ;
        RECT 61.570 51.375 87.310 51.530 ;
        RECT 62.355 51.230 86.525 51.375 ;
        RECT 63.140 51.095 85.740 51.230 ;
        RECT 63.925 50.970 84.955 51.095 ;
        RECT 64.710 50.855 84.170 50.970 ;
        RECT 65.500 50.750 83.380 50.855 ;
        RECT 66.290 50.655 82.590 50.750 ;
        RECT 67.085 50.570 81.795 50.655 ;
        RECT 67.875 50.495 81.005 50.570 ;
        RECT 68.670 50.435 80.210 50.495 ;
        RECT 69.465 50.380 79.415 50.435 ;
        RECT 70.260 50.335 78.620 50.380 ;
        RECT 71.055 50.300 77.825 50.335 ;
        RECT 71.850 50.275 77.030 50.300 ;
        RECT 72.645 50.260 76.235 50.275 ;
        RECT 73.440 50.250 75.435 50.260 ;
      LAYER met3 ;
        RECT 70.170 223.665 70.590 224.265 ;
        RECT 72.930 223.665 73.350 224.265 ;
        RECT 75.690 223.665 76.110 224.265 ;
        RECT 76.080 221.360 76.660 221.370 ;
        RECT 74.660 219.400 75.160 220.000 ;
        RECT 45.770 218.030 46.460 218.730 ;
        RECT 75.920 217.050 76.920 221.360 ;
        RECT 3.120 216.050 76.920 217.050 ;
        RECT 3.240 216.040 4.340 216.050 ;
        RECT 44.290 215.430 45.140 215.750 ;
        RECT 44.410 215.420 45.060 215.430 ;
        RECT 36.510 214.660 37.110 215.210 ;
      LAYER met3 ;
        RECT 37.570 208.130 52.130 215.020 ;
        RECT 25.470 133.050 32.360 147.610 ;
        RECT 34.210 143.850 41.100 158.410 ;
        RECT 46.330 153.520 53.220 168.080 ;
        RECT 60.750 159.180 67.640 173.740 ;
        RECT 76.200 160.340 83.090 174.900 ;
        RECT 91.310 156.890 98.200 171.450 ;
      LAYER met3 ;
        RECT 66.380 148.410 84.060 150.620 ;
      LAYER met3 ;
        RECT 104.740 149.140 111.630 163.700 ;
      LAYER met3 ;
        RECT 64.170 146.200 84.060 148.410 ;
        RECT 59.750 141.780 88.480 146.200 ;
        RECT 57.540 132.940 90.690 141.780 ;
      LAYER met3 ;
        RECT 115.280 137.780 122.170 152.340 ;
        RECT 20.910 116.240 27.800 130.800 ;
      LAYER met3 ;
        RECT 57.540 130.730 64.170 132.940 ;
        RECT 57.540 128.520 61.960 130.730 ;
        RECT 59.750 126.310 61.960 128.520 ;
        RECT 70.800 126.310 77.430 132.940 ;
        RECT 84.060 130.730 90.690 132.940 ;
        RECT 86.270 128.520 90.690 130.730 ;
        RECT 86.270 126.310 88.480 128.520 ;
        RECT 59.750 124.100 64.170 126.310 ;
        RECT 68.590 124.100 79.640 126.310 ;
        RECT 84.060 124.100 88.480 126.310 ;
        RECT 59.750 121.890 73.010 124.100 ;
        RECT 75.220 121.890 86.270 124.100 ;
      LAYER met3 ;
        RECT 122.350 122.410 129.240 136.970 ;
      LAYER met3 ;
        RECT 64.170 119.680 70.800 121.890 ;
        RECT 77.430 119.680 86.270 121.890 ;
        RECT 31.810 115.045 33.410 116.595 ;
        RECT 66.380 115.260 81.850 119.680 ;
        RECT 0.530 114.410 2.770 114.870 ;
        RECT 7.470 114.410 9.070 114.435 ;
        RECT 0.530 112.910 9.070 114.410 ;
        RECT 0.530 112.330 2.770 112.910 ;
        RECT 7.470 112.885 9.070 112.910 ;
      LAYER met3 ;
        RECT 16.910 99.740 23.800 114.300 ;
      LAYER met3 ;
        RECT 53.120 113.050 59.750 115.260 ;
        RECT 66.380 113.050 68.590 115.260 ;
        RECT 70.800 113.050 73.010 115.260 ;
        RECT 75.220 113.050 77.430 115.260 ;
        RECT 79.640 113.050 81.850 115.260 ;
        RECT 88.480 113.050 95.110 115.260 ;
        RECT 50.910 108.630 61.960 113.050 ;
        RECT 86.270 108.630 97.320 113.050 ;
        RECT 53.120 106.420 66.380 108.630 ;
        RECT 81.850 106.420 95.110 108.630 ;
        RECT 59.750 104.210 68.590 106.420 ;
        RECT 79.640 104.210 88.480 106.420 ;
      LAYER met3 ;
        RECT 126.320 105.490 133.210 120.050 ;
      LAYER met3 ;
        RECT 64.170 102.000 73.010 104.210 ;
        RECT 75.220 102.000 84.060 104.210 ;
        RECT 68.590 97.580 79.640 102.000 ;
      LAYER met3 ;
        RECT 22.320 82.930 29.210 97.490 ;
      LAYER met3 ;
        RECT 64.170 95.370 73.010 97.580 ;
        RECT 75.220 95.370 84.060 97.580 ;
        RECT 53.120 93.160 68.590 95.370 ;
        RECT 79.640 93.160 97.320 95.370 ;
        RECT 50.910 90.950 64.170 93.160 ;
        RECT 84.060 90.950 97.320 93.160 ;
        RECT 50.910 88.740 59.750 90.950 ;
        RECT 88.480 88.740 97.320 90.950 ;
        RECT 50.910 86.530 57.540 88.740 ;
        RECT 90.690 86.530 97.320 88.740 ;
      LAYER met3 ;
        RECT 31.560 70.810 38.450 85.370 ;
      LAYER met3 ;
        RECT 53.120 84.320 55.330 86.530 ;
        RECT 92.900 84.320 95.110 86.530 ;
      LAYER met3 ;
        RECT 43.670 61.140 50.560 75.700 ;
        RECT 58.100 55.480 64.990 70.040 ;
        RECT 73.550 54.320 80.440 68.880 ;
        RECT 88.660 57.770 95.550 72.330 ;
        RECT 102.090 65.520 108.980 80.080 ;
        RECT 112.630 75.380 119.520 89.940 ;
        RECT 122.070 88.300 128.960 102.860 ;
      LAYER met4 ;
        RECT 70.230 224.095 70.530 224.760 ;
        RECT 72.990 224.095 73.290 224.760 ;
        RECT 75.750 224.095 76.050 224.760 ;
        RECT 70.215 223.685 70.545 224.095 ;
        RECT 72.975 223.685 73.305 224.095 ;
        RECT 75.735 223.685 76.065 224.095 ;
        RECT 1.000 222.050 45.850 223.050 ;
        RECT 78.510 222.110 78.810 224.760 ;
        RECT 1.000 220.760 2.500 222.050 ;
        RECT 36.735 215.190 37.085 222.050 ;
        RECT 44.850 218.650 45.850 222.050 ;
        RECT 74.770 221.810 78.810 222.110 ;
        RECT 74.770 220.000 75.070 221.810 ;
        RECT 74.660 219.400 75.160 220.000 ;
        RECT 44.850 218.140 46.390 218.650 ;
        RECT 45.850 218.110 46.390 218.140 ;
        RECT 74.770 217.570 75.070 219.400 ;
        RECT 44.530 217.270 75.070 217.570 ;
        RECT 44.530 215.755 44.830 217.270 ;
        RECT 44.335 215.425 45.095 215.755 ;
        RECT 36.555 214.685 37.085 215.190 ;
        RECT 36.555 214.680 37.065 214.685 ;
        RECT 66.380 148.410 84.060 150.620 ;
        RECT 64.170 146.200 84.060 148.410 ;
        RECT 59.750 141.780 88.480 146.200 ;
        RECT 57.540 132.940 90.690 141.780 ;
        RECT 57.540 130.730 64.170 132.940 ;
        RECT 57.540 128.520 61.960 130.730 ;
        RECT 59.750 126.310 61.960 128.520 ;
        RECT 70.800 126.310 77.430 132.940 ;
        RECT 84.060 130.730 90.690 132.940 ;
        RECT 86.270 128.520 90.690 130.730 ;
        RECT 86.270 126.310 88.480 128.520 ;
        RECT 59.750 124.100 64.170 126.310 ;
        RECT 68.590 124.100 79.640 126.310 ;
        RECT 84.060 124.100 88.480 126.310 ;
        RECT 59.750 121.890 73.010 124.100 ;
        RECT 75.220 121.890 86.270 124.100 ;
        RECT 64.170 119.680 70.800 121.890 ;
        RECT 77.430 119.680 86.270 121.890 ;
        RECT 31.855 116.570 33.365 116.575 ;
        RECT 6.500 115.070 33.365 116.570 ;
        RECT 66.380 115.260 81.850 119.680 ;
        RECT 31.855 115.065 33.365 115.070 ;
        RECT 0.575 112.325 1.000 114.875 ;
        RECT 2.500 112.325 2.690 114.875 ;
        RECT 53.120 113.050 59.750 115.260 ;
        RECT 66.380 113.050 68.590 115.260 ;
        RECT 70.800 113.050 73.010 115.260 ;
        RECT 75.220 113.050 77.430 115.260 ;
        RECT 79.640 113.050 81.850 115.260 ;
        RECT 88.480 113.050 95.110 115.260 ;
        RECT 50.910 108.630 61.960 113.050 ;
        RECT 86.270 108.630 97.320 113.050 ;
        RECT 53.120 106.420 66.380 108.630 ;
        RECT 81.850 106.420 95.110 108.630 ;
        RECT 59.750 104.210 68.590 106.420 ;
        RECT 79.640 104.210 88.480 106.420 ;
        RECT 64.170 102.000 73.010 104.210 ;
        RECT 75.220 102.000 84.060 104.210 ;
        RECT 68.590 97.580 79.640 102.000 ;
        RECT 64.170 95.370 73.010 97.580 ;
        RECT 75.220 95.370 84.060 97.580 ;
        RECT 53.120 93.160 68.590 95.370 ;
        RECT 79.640 93.160 97.320 95.370 ;
        RECT 50.910 90.950 64.170 93.160 ;
        RECT 84.060 90.950 97.320 93.160 ;
        RECT 50.910 88.740 59.750 90.950 ;
        RECT 88.480 88.740 97.320 90.950 ;
        RECT 50.910 86.530 57.540 88.740 ;
        RECT 90.690 86.530 97.320 88.740 ;
        RECT 53.120 84.320 55.330 86.530 ;
        RECT 92.900 84.320 95.110 86.530 ;
  END
END tt_um_oscillating_bones
END LIBRARY

